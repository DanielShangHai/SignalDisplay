t-�'�ij��l�˨�w����iKHz	���O�E�qM�Pp���%vE��&Sv;��O-2�}z�fgX�w�~[�����쉊:�:h�Mo�h��A˴i�A���F�l�����|aF`>�#��T�*7�¥�����s�q�O�@��.��;��4ew{M�� _�|q��m�Vr�W��!w),Z>U�̋�4oa�|��v$�,E��)C�����%��Rn�� /|�Q��9�l��.����x#�����IYlV�v�s�$BQX'^ ���'[����Ţ2�B4�����6�
�n��p����N��ߐ�U�o8��c�ǳ(Ӌ��g��z�Q(�3m{1��;��_r���} ���	ұ@��������{�+��}es3q������}�/����R��/�y�����7�lT�c���dA1�哣��Z56�VSxg�	�������hilQUæ�-hI�]>2���c��_�DY|H�EC
=��`%|��r�B,��L��fN�MNR��1�a��ۘ���l�����n��|�]Y|ID��A��G�@��d9����S�|4�V��T�$qNB4	�-�-�2�[��	Qc�N���r����d�����-?��VO���0�C2NV�x-IL�N2�͋E�9�J�jP��d�w��
������z)VL/J�GM�Ԧ4^	��òX����4��h'�^ZkL�HֶW�	
{'a���:�]�yD��?�T��(x�D
�9W^�T�-�rx�V��82��DYu]����@{�����Cۙ�6�碨���`Ax+:<tN	��1X�t~�2|��P�xD^��ۄ�����k�P9p~
4H��|�['�-���h��{���(��[���VX��������0�
1�u�L���E�UyN3����(��'ms/�)�ܚt�Vcm��h*pFw��B�hH��M�{��e��C�[(u;V{�ab
��:������	�������Y�_������|Ư5?�b� �mwK�	J�s�8��3�����!�T����a������	<��N�H��������91��x���ݿ��Y������e��:W��$��Β�O.n����1["_�F�.x`�M��l�Y)��Z�Ķ:��,(����|u�Y����٪�A29�/��_�$ (���/��&���X|�~3ߴ�����mv[�/�4���GLpٖB��jz�����D�R�	q�F�'v��[z̬�W�IG��4Sf�)kPXG����+$w�a���r��-������:"�3�J��D<�l	�|2�<@R8�#_lyX�D ��O>(�ms�6v�vFM��;�nD:�����H-$G�e1�dL�G'�����f��@��������P�e�g�;i�сo�Y����3�}��Ύ튓	~�
D��:+D-;�Ui���HC��w�7aq�AcV��D�Ϝ���HΖ���^��	/�r��3:L�=�~��G�J�9yzz�I��\�'��t��^����������ɑ�nR�| ��&G��WpR%�c�U��q�:4-�\�GK-�7��	G�����0��h�eb�Hht�g������w#z��P���,f��6�?�g//ʑQ`� ����ϰ2���ӌ{�H�B\wX�X�o�P="�+Ʃ��6��Ԍ��
\T�1`��=��ݗ�Ji0Dm�o���ceC`~ �(����t�e��Gς�yr+1F�X��(x����>�n`@|�c����`܏��&�Ȍ�����~́[��6�_uU��,<�t��"h;z�a���S�:KA� �8���I���͇�|��$wa������m���taD���ŉĮ!<�5<ʶRE���%4%���������8[�GQLL����`�K9��M���s�'r�H<�P��	�#����a�����`�f��h>������C��_�t�$��mYa����z
^�=��8���H���)���(�$�~f�>
��P	˭�BςRd�ٷ96EBO�{�a�o��e���=�s��~���a0�9�>)/hi��� ��-���������tz�/�k���+`o2�+C��Qtn��Z�/�;���ϓ��ؐ�).Ǐ��H6�5�Jݔ�O�j��A)�r����|�y����k�Zw�Ԃ#�V��?*S��)'f?�D�D�`���A(�� z�,�o�ݵ������p��Eh�jDxf���[�������y}��h�D5[�����r����J#�@rI�E���;�m}��Gf:*l��jj�����	FFHF�k�
�s�g*�n�S6|hn����rw�Ks�v�:�[w����|��ۛ�&PE�?����ڄ��I�W�!\`���CM��������0��g
���6`To6� >�=��e��F>\dAH�H����"��Н���^�g�r�����+��_����)����Qp:��Qc��gد��<"v�4���n�@��&�X�A��5,VhD4x4�������z��a�B-���X<Ӛ�� H�F|gЎ6�pZ3k�|��M�E�<��;�a8>�]�2�L�<.v�r;�R���H5�����a0V�@�
�$�AM�I#�c���$
��o�&�}v1�F ���&�~efw�/�$�צ����aeg�,.���ȉ�zeE@����i�7<��Am�p�fW	���>!ς��|���¯�+�;���+�'JC,��}l�{*K஠��D�@�Ԕ�.����н�!}��k<HC�f4f�������f�抦�-�{��.��L�o �
m6�U�	Bٝf���A�ϫ ����jj_m�?��R��9�1bO���t�v3*w/�ɻF�S=���X��zd:��|1۹kh
��BX$<m�c÷@��k�H��셕���$�=/���a�vC�-���t�aJvмAY����zv�XY.hAe9J鿂}��M+O�**A��pn2��Dq����3���Ln��[qUL��X!�2D�&�·3M�<�_)ǉ(P�V��/|<q	���i�gD��Fu�>>g�a��:�9����g�?�\�ET=)WK�3��@�܏�_��mi��A�!40UK�/��:e:��hL�+�e4�.�BAFN����l'e����s���N
�%g��?Ƕ�$m�C)���pD"_�C,��Hq�m�E���VF����g.<�R��:�;��x�ǃ���|b_c�d�YN||�VR����R����V��)��:��$��
ଭ��n�G���"f��R�f�w��b0�2~��D�i�>s�i��3��1VW�M͈�os��˖��,E�M�4��5L@�ڮA����夆��-�E=p�{̦/��33�;/z��!ݏ��D�a=�
��Tk���`�q����;������2�7�0��,}Sɚ-E�u�G���.�������b	<���\pk�Ot��& �">�~��HS*���0��!q��8Aՠ��xp��ݱ�c��Kf��
��9&��l*cO�;�(S�r���/��B�{Q�o@�-�3��/�A ����I�nq�8��[� ���±�G�
:V>bFFS%�YiG1�i*?^\*�e̦2�}|���f��@���}ʤ����8�dd۫OZG��D���h�0vD��/�!��߿@�r����C�E|X���><0�ȶcME9�����������vCX�w๟h��i���7Ivt���jb�g>	͸ie�F�
�TM2ϝJ�	!:W�L�ڟ%��g�_�3J cx��CZ/�?z-����!T#P��_�S���g�	��d�/}7�\�[Ҭ�ҹ�V�+_
H K�ջ$iV��ұ���2_�%��!�&��(m?�j��1d�7�@����4=S�_������0���#��}�"!	�"T�?�]E?r����qYq��e��Ċ;:Ơ���� ���Hށ�/��cp�x�\�॰�Xƶ�U�����s�*(��ut�#;��\���v�!�������Q��}o���G �'�ވ���3��c�ƫס�!���K�D�;�� �2���l�JCk��#G������<��|��(�����W�!,c�O1\:T
x6�H�}�ԮHW����1�l�뉿�	-���ˉ~�o��m1�N/%�y�4���8�50Jv_I���˛AAs�ç֚A�]�)gѰ�m�$M����w�)X<J<�}V���-T��f �0ܰL4�1�O6gW��[G2�C$4Z��q"���e�	�ڟ��N��v�ޒ����7jz���t�f��ƂR��C�n?i������$��7N�*z~2���5�\դ���b�M'j3��yD���R�0^�>��P�ug=����@t��Í�7ia��1�)������b�#> ���G��hU�h"(����B��D��6z
[�0nܤRm��$Z�	.�s�"1f��+���������p@	Y0�}ٚ���.B>�m:6�g��x}��Wx̓�	��c��_z�kzJ�T(�f�s9�`T#��K�݌l�*�	���2_�b�$�/`��:M&6_h�w�LEM+���</,�m��Ï][ҦpU���k(��4�:�z˔�r�:Y���pJ
���O�w���!����tu���]�߅��Y�+�eA��M���bo��O�����$��f_D��-�Ƃ���ɷ��b+�\A�I�ݟ^2�z�p$i^-�R�$-�(���i1�m����ݮ�Y�������9=����F7��釤qZ��Jj�3�x���$ʑ����&{w	'v�>߸P�Pdtv��&��-=�|Շ���*7�Z�˔�:��d�M��]�����W��vf���E>۞���c�bR0w��w<�����������,$�a����5&k�<;�O9�RQ�� �Y��B��	9�@Rgd��3L�����(7l<}�;	x�U�̦�0�Hi��\���%�`㥧$�0�zi@�˾�(QV@"g���C���n�S�~�%���g���M��44\��p�-�e=@���x`��,X��-��<9����	�m��<ֶFD��;��#�����ʆcl@k^寇�A曀��#B@�ɽ�Ӑ�H������f�F2YÙo��OL�Ix ��=C*r��g�dc�[ˉt�J�_dlc"��0�d4�M S��IVs8��L5
۶��Q`�@�W�Q�z�����X4�m�͗�F(Pчne�D��5K< ʶB`�y�>#����$���ʃ�~�2r���J@$��3, 9����� ;�3��1[qw&���/���
�
�;���iY�S�҈swy�F�����&PHs�|�:k�1m�:��*�Z`��Jwov�;��T	�hi1��_I�D�P$4�Պ��'�����>	3p(-,�B��}ْ�Z��|*u,Ye�Uſ�L��8���-����J�A�Ӷ��ʸVb��(f,ȁ�{�j�T�F>-�v�"�Rs�jɟa࠘h���a�U!��e��	FMU�9�����g�8��j�cϸ\e�S�7*�_e������b�=Z��u48�#&B{��x�Spl&�%��3D�z�����yz�$�P��ɣ����(ip�ny�[�4ͼ"�j b�6���W����e�',�c4r���o�EO�4�4�$K�����O�0*qꢒ�\����)O��c��1�%*�(�A��n{�~\p�!�����J^�A;��d�9T��P�Aؕ�?��Q0W7�Z,6=n������q�g�X�r�`�1S,;���_wr�	�/P7z
�6�*���@�>
���PsP��f��(��ӯ/������.��~?-J���7���������ӝ#��IV��߂H��TU��_�U?1���0z���T�����6�>f.�;����r��(���7��i��9�e�pP�g�����xCޡO�&Wi�.78C/o7�PڨI�(jqoœ:�4�N���@�
��ؠ. 6.������a�e!��4t W�S0(õB^W�<(C�}�@{F�*������@̽�|�&��4�^l�@lW�y��=���G����Q�Aȑ���'X�j>��1�zD�D�L1�"����dÐcW��,"�oB
���56��ڢ�E5+a�3��F�u2Q7�I�d��%T�w��f���5=�	ް6*xQ0n��z	=�o�g�2�9P@�:*�-���mq�ȍ'=)�3��V/
mƩ!=��e6�;���,8x�mN�+M]�3��pX����3]�P��ۣ(&@d�_�|�l���&`�2R�1izW�er�@�A�Y�8Ω��پ��DH���u%��kA�Ã�C��щ{��I�JM	 *@m�Dt<��֛�2)~*ݟ�G��u;0R&0T�P�������e  |ca� �!�!X�Ns[��_ǝy�a��֪�ь���~��a���߂||�@��4 &lF̿ݸ�=@������#����� ���T����LM��.�@�M'���+A�f+�͕�$)�*�F4�i�4�F�<�}."<.�$CɊ<�?�,v⡅C������cмD�m���#�w�ȥ
��݄�Ec�Lho�-���������p�׶n������������^�ll:#���Ne�
\���A�&2��/�P���U���������d`�REx#�����mW��T�	�P=:��l��8�BR�A�?�����~s�{N����Lk�����q���Ŧ�D�9/Y r"�!�p�L�e�D�ER�ʀ�%V��&�����#"d�?��1�{� �� ��F���U\�U��J�%l�Gzx<^�a�4�l�QS���
�4L�!X�~����2D�ڛ��<{����V�c$lF�0VWvZa%�oc\d`��Ř�sLYDrXP����1
#!=�vxq�X������R���wO�܎��!j�݂�B����0�Cu���z�B�=��#���6!�?���:S�g���*��`p��� ��������$�}������c��#��BL%�PI�'Õ�C�������el�	ds<����N��a�.�릙Ail�r����h�w*[����W�O������ 3?���x�э5�BT6F^�#�F6:�%;�e�)�8�OP��k<\'��p�%_fD��	}M�젦7���n`�툘X�F(c��Gel���7�>�M��ZZ��*E��"J�_�E3v�&`Տ���A��Q�rż�a���v�G�޵3��G�����LS_3_a;�OCf�Rҡ!�J:e׌�k}�����m!�5h~Շ��s���֝?�G"��}�6 �Z��5��Sh�P,5�U"��Z׮��cVvd��	� 1��.�Zn�n�.�������[rn{���PYږ�/
V������W�	|��![iQ�b=�ݙ�u������=��s[=-Q:f���/+���µo�>_b,�ȓOO"F�t}@{.���Q��"LN�wa���7�V�
���]pm�{�N��WpBVN��Б�$�Խӓ�5�5"��v�:�M��������x�<Q��@��7��<8�7��k�biG��
s��=/���0^��;����!2O�h�n�UC�����o��i���\��P��c�!g�`S�d��޾��")��|�U���r���T��Q|�2�����Y����:��pF//;/���Djs����_�jO�Y��7���M�9MY
U�����3a��a��e�|`�aN�𢪽���>P\�d�/���,���Q�����aX�^�̋��ӌ���)
v��_k�xò��bMt��k��g��;�� �7LG͙�2���D�(��ǰG� Ҧbz</�T�ɲ��Z��.# �m<��'����%��M�
X$xoBl��^��ȉ����*<u�eI�^�<��4�eF�z.XLN�{F�S����D; ��:�̩>�YB̊�)���7�O����$�J����y��A�z{���{�@3��	��{�a�����˻*I�XqYt��pIm�H��V{ώr�q6V-��!_��c!��A�K�����&XhD���tŜ��a)Z�|'��FJ�
>���3a�o��u cr���9Xd!�5�ONr#7y�f_Áq���:�6�����R�����s�5.�䇈��,(m�����dl/�ā������}Q�.�ۑ��u�+�1'���
�!C���\�_qÃ?���b�}��7�-dΌ���U ~��,aAY\��%�k-���J `^%H�������A��`x'T�n
S
8���b��	1]�W�9U����� {�C���n�8h&t��.��.�R�`�[@�r���I�)�G)N`�G�'��c�}�]4e�N(��_|�>/ľ�(Pf��g�����H����XxH�0A�~ϛě��*��r�2G�>��������`�[�P`�@�`��<�.�vNe�~Z���zQYM��wr�D-���Bzy|�i��H��T��'9���Ї��B�X��l��uZ���n]SH�Xi8�d�w�48��=t���n� k���!�kZ4���kj�o�'S�ُ�į�����(�Ї�N6�e�P�����mo������6�F|����ޖ���	[���8���fhj��Qd6:��(���V@�B�k�x�H�RG#�/�Q���c<S�܇S��j��c�¦z���M]Њ{���ɯ�~x�K�RP� ��Yq�!}�5�祈��OOϳ���4�v晍���_�GcW鱂B����H�� f��hb��{���h)�c�:G�Nl�6Z���U�s_`Ht�|#��J�
��[^�$6"|# k�Q#&} �ҬDv>C���Z���2$��a2��:�D�4m_����6�0k�v/��mj�`Q�p>���,���}�J�6�Ob�بc�S�� ��iŬN�Ek(���sM�uq�_�7D���XH�T+��1�'��(e�*o����� `��Q u?�/���F�ap�`�M7� V?�P�%-�Oa~�y6Jab����&U��~��*GPL���q��v{ꤗ��� 4h'��o[}����n���f���/v1c�F��ܻ�3yG��<b/j�;��D�<(d����w���	�/ �x�z�z�[n��*� �HHl0
P+��%�fvz`���O
�e�ہ���P�*O���
�!@4����ި@*��i��*JF��)_��T2�I��V�R�(����C��W����
F��E���T0�'Q9�G���W�	P�wz��;Ш�	�5}��;��Jr	;�92<bU���?���s��#vL�סN=�~�B��DU&]�!v���e��V�m��{�r=��"%*O����}ٰ�3Q�A����ak��6R>sp��+�;�_,: 6(�DC{�PJ��Yb����1ĢB�e[���LR4Jh�NaT:��&�t���PZ�j&�`�j��@���jy��n��>b�3��2�s�ƅ��v�Ze�)Ō�D���[N�!!a^���'���eA <���1��MW��sY[���DXPG^�Ѯ6s[��'���4�n�@�zh��*Ǡ��\���4\|@|��?��GG��l?L~��8*�`�c:��??��
=�.�hz)e/�E)�pp��t�R<p�!�c<pԷ�ߌe5s"���%�7}JZ���6~_!�c�.��=��f;���ဈY+
��Q��nOP��uVy6�+������X�_GX&+PvJ��p"���`�" �>2;��y>��Y�d>9l�j���k�! ��pm��~_���C"P��GG�� Bhҭ�p��ћ���Z6�@>��
�J-��1��	n������7�?�ч�����ǌ��t3�1�G�Lo��;^ *��}���x`PT�Z�ۆRŗ�AbI�����s��p���H4�����}i��l*��<T���И��($����yq/���2��c�q�I����s�{�r7pF!����	�-�h����a��.VS����(�R�:�j2ܿs�L
�d�p�KZ�Mx����Œ5x#8�ݓzA�5)=��E�@��I�ӈ4�nwikN�X�z���yf-�'�Ĝz�"1�柶��K�vF�>���W$�OH�0�EA �x:+��0�� j���>�_��(���Trz)u6���9a�n=����uE�� =k����!�15ci��ȴi�>YD�}�q��*h���-�kg?��e��:��m�ؘ����9���Z��#c����e�		�@cU٢+
��dN��KXvH��腕�+{)}�F�m�����G�
D
�,m��JlM�=�s�n�$O�ѡ����SC#��/��(�"k�I��W��'�	�әj��N,JD<l]��csё[�bQ;�t��^UE���"�G�ǐ���0d2PN������͟����._S�8`�9�*�Ǯ]���|2�~�("g��%f�<�9���gZ�����|��._��Y|��D��_!DR;_G{i^�A �
�Z����ȥ���=�����Kuk��Ƌ�b�YW���ݧ��!L�|�Oa���%��U����P�2"�1.����0w���ɕ��4�	�4���ӎJa��` )|JݱJR� ���GYf�yЁ���j,2����TC����#?.���L@9�W�DƆ�]!��D�9��@
�np�ji��\�%
k�Z�(��*��T���V��g�� ��a>�q�;N�-&���R1�z3��ȕF�Ap���P�	G"a@�HfA���)�r����G��P�gcC�ك��f�9�6e�'H�3�t!y� 0f�7�Txq���~����^��h�$ۉy8@�N�.���ޫG�~���^�?����e��dVQP���S;�4w��*����iN#�()�=�ݧ�r�xa��͌��!��M⃸L�c����B��i��2)��A ���L	XeNs~_+h��z�gڠ�����!CvR���l�S�=~���h]&+/��z-��'T�͏�}��j���T���	'� �̯$��8x�M2��uQ�EK���� ��А�{�<�t`�W�r�Uз�!n�kB)�X$,�J�U�����e����"�+�t+�_'�IF�t'�Di������������?)#�	w���������I�Zp�^c�g�� m�7
���7����X�Jd�-��������4�x���6�!�,��T�yd+���O�#C�oCG,)�*��B,�~]UV
�T+���*<m���B����\IE��-�/E-�>D!dж��̏#�W�@��.D��,��?���q�I�t�\���JX!�O�\���� �L�B�+k�E��/�֑Z�f��
R��M��=�a���f����6�'	}#4�L)�}͝񂡊� ��U��u.�)��AX��}�0�+�U��UH�O4�bB��/�ԍ�%��U2�d�X��(Ys/k���DK��|���(��5�
���r�9E�}�Sl�'����>��$����*#�\�آ�y�?�'��-���t�����"�k����c�|�_��L~B2"��D�Ľ����sLt��{)�	;G/��c�N�bNd�;�����N�=����M�e(�C����p��|�y%��Zɵh�%�ߴ�'/�KnFU>>����3-�0��x$��f=�g����ܴ�3}s����Ј����d��Wd�*k��J�
8�St���.���M��>��*)i�M�Wİ�q��I�Gz�I�o� �i�(Tk������a+=�5����`�%�K���='�ký��b��B���ǎ�hq��0���3�p!��aA�%�x?C|��t�&	W�
�7�[�,���/B>��O,t6�Ҍ�����C_8�Sc=�1(��nv?j���� Qn;ș�H�wBD���!B���Iw�q4��e;�����-��i��?r�՝H�m�4��ؕ��l��X����D��B��
���
�������<�dS��M�}��2�ϑ���2�Rs�ww�B�	��!�-��Yi���{�\���v1����n|E�
*m�X"�[�]� ����Ee�������?^؁(��#r'U��s���Y�����XH5xV���"���A	�L��b>����K��� ��3D_a�K��!T��f��(B�����N�+�:9?XDa
{�ڦ���\т�)0���R�#�u>5��=f_|��#7rf�r��k�o,Z��%y5�\��pN��Wv>�>����N陾v�����(�AEcX�*_EN|�;�֑�D�v���&��F�}��I��o��J���%H�!�������0T;K�K��'ǭ/um�l$#��E%~U\H�3���0��!t�w��3r�r3v� |��1�;ؼɱ�/�;38��*�A�<�����) L1�?E�~Po�����m,�{o�jn{�{�!�$巤4p��ӷ�G�>p��$��࢖�urA;�*R ������!(@P���!=V~�)�C��8P)�K�)��D�[L�E�LW�.���� o�aV�E罿�:�2�tD�����X�Ed@��Y���8q�GTfT��V�@[�fkf�j��?eC����++"w�Yp��U�#��|!9�R��j44%
	
��!�%�		�C�w\F[~$���Caĕ�o�fJ��X@)1�a��p�Θ@�a�1��wU!��7�S� ����!��J\��&q-�8�(??܌[��1\@�~�/l6c������8���[� HaD>��z=�N}�Vⷊ֨c��a�q:�R	��a��?�B�e�q�$A�H4�-���֤����C����s�6�.�_N�0�)O�R�����	��T�e�\��ţ�������|;r�8�yhC�(>n?N�_�+)~�����_�������D@�ق	�@eA�\ ���g�S6����r��71j��S��eEJ�!�2%nY�}받���=B@�Z^��a�5�t�o<?�m�ܐ�XP����Ua��r�����}���,�����t�tQ|�ѷ��"o�L�Q�?`H1�_IM_��!Y�！`"��2�קԷ��c4�3C�@��Aș��쮾�x�kH�)��~��$�
v��8�l	,*D\ *��i��i�ɓ+j3���p�vf�� ;{��0{���-��|��TW�(;NjS㽴p��T!�¹5ڗ$��iY��M��`�C����$c[{��
��Dه�AJ'A�XL��KrC�v�R�>^���Ŵ���(��U U�	��U�a���]�����V�D��5H��/�R������i�Ӡ���Nx�>�&f��.$������� HO�#�����E�?z�ά�_�Y�MB���EX�D���x���φq^��ꚑ�zQ��O���j��Ag��>w�쉥K�H��^��_ J�n���r�\���o�3~�K
��}
��ŵ�`��NO����Q%��ҳ_W�}�:+%�X��t�0N�O��?�{�l7��%=���Ɔ�T/�-�O�/P��XD2Q��E�Tc
�Pr��v���_���8��/�q�0x�̓���we����/ԥb�ന`�J�����8����3�� ����&��x>Y;z���V8P�A}�;��8�-/���9׎�7i��X}����r1�`�Sy{o�r��<�V(�Q�����Ԃ�p����Yג=oQ���F���%���t��[��#}�?��Ķc1"xF_�!�1A��ϣX�N�?�Q?�1m���0��ۑ���r������o�]�_.!	(�G���\ӵ�
�RF�l8��-mI��a�f����c)����Z�y`�P��H�}-���#a.;�_�'�5>�XO/��p�`X{�y��;��yy܉�#L���È
	�"���/�R���z�iyHi<�0@�AR�(s0��zW��R����>�<H_~�XصAQ�G;��
����E5��Q����*9B��^�A�/e�D�	��<�X���K�@�������Q��wu�J_bRy�}�����Ц_.Q��s�&��0��p�M6Uv�<���U�X��\�v�O�/�lJ&Ԉ(,+�	FN�WS���;mgM'a""Î�Ȉ��m�Ӌ�k��\��|gY��!hf��e�f&V<�#"߈�R{+F}�A���2LhT"�IPN(�ݐ�V6zg�,,�(�L�|��)s��/}��Eq�Xc�D��߮�Ա��tR�`��ȏ�)��� ��"f$84
+����;e󤃔����x��B�ʕ2������˓n��;&�m���+�e�ݍ�:�&��z���d��C� �\:M�u����e��̉9QAO��?��V�M�Yb^\AA�e����a�_���_�Hw P~��2���1{�=n�˃c#ųWe���|�ꄍ�sI��(W�s.�/2LJxw\���0>
���u
����wJk�߄/�ű"[wp&h�;��j%�����!,03�������j�&��7K�!`���lj�������'n����Q�t%_�*8a�*_�

�9�L�=_�Pi�*)��Q2TEy_������Q�}���j��"~hE�6�`��ܝk�Y�F��䟙oheo�LVH�a����tM���I���_���������]��?�a6���)s�����.��Ǖ���BhA�Cx�M��/��<����?|]OO�$���k+�>am?/�2`�E�D%8��ĠL�We�Q$[��HQG�OM��e�r�N�!�?����%�&K��ŗ�-#	���r	T��cn>��
p�����{���#� PH��pn�?�����,CE �?!��x:�a�,�h����6�$_
���%`y�l��p1Yh�q�s�&ty|�	^n�l2*�G��+ cthF4o�MҢ��!�R[�K򩄳��� ]�R���`��E��
*�?n�Y~��J��Zd�ҩ}�_�!�"��p�֑ �c��i��:&�B����W;}|��F4�A&�G�|�!�Bhڦ)p���M�(:b���0�8�>�s_�7�,,���3��mu����h�`��?@������&ۛ�@$�{��Q�W���?"�e��Ke�))]��:�2���l��3�܌�~��`ߠ����믩[��1q�w��ʿN���-���^���	�7�#�rʾ����=3�ZlVX^����N_/\�o��PH+����/U���\��N�����7u����^+���,���9��S�j0��ۧ�3KE�	�M.�{��پD�W�eT�.Df�s��2�o/(`r��3�ZZ��QT�഻C��I� ��C�� ����)���;���8���1���"���M�&9`4��[(J�M�{N��bs�ڴ�F%n� �Q��a������}��G0�		|
�T�Z���N��T8��T \���Ba� @����f
��}��\5�aT�V����/��P��-��!�B���AǕ�B0k�/���પ�V�XfH���Vܥ�0ʙ��X0����"�z�9El��쪥
�Ga錨�$��N�b��+���j�K,���/�sLbS#Jd��r��0���7󿐁.��BHT��	I��i��H�p��Q%D�$xw���m�׿�!��U�TAC+�F�6��3��9���p%w�m�liE70��[�����=|!f��#�N-��'�Z���]6q!5-�8$q�&?��\(B4:�54����̊�-[�BL!� �f[E��E�\t x���s���DK��o_��~'��!!3n�z�;�"K���_LU�;}˙zw�L��e�	x�'cX����T���?kavx�%R��ra�b��_��%��+R�g���ڟ랦I����s�\�o�Nk����q܊��,�`�:�q�!/���?��+�|�E	�2Y��R��V����~&���f8!!Df�e�EZJ�z[@v�F"dC�K�b�ŷ5���}_/�9����q2@8�^�����>OtN20�oe)|AJ@�l�A)e�}��ۊ��
X$}C�lXH�`����;-�S3C����QB�2��	��r���f��0Ñ@���/1+<n�q?��8����|S �� ��W�l���զ[:�6#qOK�t�vٺ8e�,��I��ɂ�r�8�*=T�M�Ku%�<$v�B7��x���e�D&����l�P�}!x���sfʅ���*Q� u莂?YU���&wQ�`�
�!+��F)��N��S�T�h�,	�S��3�Ƕ��Lr��������{�f���1�#�y��{�"�r_�]�FZ�zc��cB."���r^�&�;�h�4K�VB�	���IL��8���\�P���a��*N���&LeN�W�|�#���
6&(Ia�hG����X���v���sS���EÉ?���g�Y�[���e����V��[����� a�|��QGqg����=��Ĝ9ܸ5C��H�*@��鶂��/���2���Bф�9�=�Q�ߦO��1�p1��X_�����Ƌc0����� �r���&����9������	��U���)A0�n�M�[��"��zE����}�)Ϗ��L����Ⱦ$̏�e��!$4M��ܢ�=��#�����q|�]�V�-�޷M��?�.^:c�⥬O�8l�6����XU��9��Hkf�%I>�D8;o�chH=(g�5x���!�q7�g�����5�r����}��$&\t�ĶG��,/�)Ļ���e��楻	ގ$px�d�|� B��A\��-���GK��/�+rۙ*\�/ۻ��?�{�.�C�)Ml��-�M&����*��e���P��O�� QA��m�F����I/0&�@�U��G�4���G�_m q�q�'���1�I�ښ��e���v���~A�&�_��h�-�Ƅݸ�(���>^u/�H��(Ϙ@��B��8���ϟ��m�yvn��֩1v\폵0����,��պϪr��K� ߸��;7��o�j��/��B8*��>0#����n3qи��B׬�`P�(���	-�W��C��b���i����s���.s�LQ�09qM�Z䴿L)ч`}i+ؼ��+�@���0��Dc{��%�?���*�x����HA��]	t�(���EC��CV~K��YOD%u9�ՠ�zB
:H\G-�/��qh���(��
�1_QL�w��JY}�I�o
|{��sd��[���K����*��i�;8t��^Lϯ��R.�۹�N���&��7wy_�H/+�oᱸ"x�T��ƥ�7��T�~ ���o?l턂NxG<#�X�Q����1�4�u]����e�̜o��0�P%�� T���c��,}����4��Dulp#j͂�aq��fjr�(�@'�鼾�$��3)H� �?��r�Vq���^��kg�0:���8�]7�d��u�gV�|��s����o/�A%��a��GV �ܬ�m(��Q����Kfٌ�K�㕍�L���傶��d��ʺ�_��T������T���0�ĩ���8������M9�_/��p����0M)�M(,�X}�#((�Mx�S����ʐ�Xl���M�	�q�q����C`�2y0���O�E�Upê�R%�,Aa���JÓ�����1��Ix�K��C����H�4�Q��|�l�F�	��y%r��D� ���M���'��6�.M��H����tz)��*�' Nr�J��Uw����0��z(�6�Lh�To/�(�bP,(Tjn?#VN\�f�|�&�wqX��w>�}�W�l��(���Ҟd�8��E���`��� ��q���q#���=}�R�BR^�~_�)�*}����G(0���/2�f���G!�	( q�	C������i�8��)f?���$�;֛�AqS�����?��R�cWi����x-´��0]�xI�s�2G��QC%�p�E/A��J �[�D#�{�d��<\5Ļ�`��J������+cC�\�^�U+oKo�{O��* �
3���KF��3���+RwX.���R�^W	E�}�PW�4R�/�I�`�������pl�Ncf ��j���5z�*�>Ӳ��M�	Tp�'V�®ʃ�Ȏ+s>5�h�*H�Q5ZG��Ԏ,.�_�J}I]r�o��s��^`�"��C���/���%��կ`�;U�?����b�I���Ǜ��A�L���/@��z�4GES�F{�C_d1JS��]���H��C�q�vc����ar�� ,�:w��_�_)r����ĝ�ݥo��s���Iw��tG����)]2<���"w�i��<7�_1]B����_tN+x�߶���+��+��o�}���L�_������z��j�.6���J��D�k�s�#����G�aN7����hh*		�M�K��wM��=�@���Vt�G���4��R�Q�@�b��<W��o��;QU|3��_4���}�vS��ZB�;v0�jKa�p!���u�������3����f3>N�C�h���a1���lvS�s�N��73\]��M���0XT ���KN� -��$�{Z�:{�vKh6|�b��M�L'\��J��������(<�Er��l�)�����(}�k	m$[�ݲcz-%8Zk���7{�G�Ԫ�@�B���I;�q��48W�RC��9���2��O0�۽���';!~��]E(��>=�ؤ<*)c^��̂��Z�c�9�i#����I�0�)B�+c�b�E� Jwl�z���2�) 8��flK�H�#AaA@�+�pۡnAf���HsA��������o�׮k�Y|&%H%�
H��K����9ݼl��{|��㠕�[q�o�6\>�xDOC��D�oŗ�1\eQ�1
u̓w� ��{[���g���Wa|��R�l�7-�0�	0� �FU�j��H�N�R��Hz.�����]��11Ҥ˯����/�8P[��5|A/k����N��ꐡ�NI�xDg��N�R��h�
��
��|��o-��6R��|*0q�PR�E��T
��!Y�:k�+<�P�w�b��z�x<lHU�X���y-�ʼ�A~�(��e�M�Q�Ah
ʬqN�x��s����ծVVv��E��yQ�uk=�TP�V_����W#�"b��~}����$M&�Vovy;��B^��ѸϦ	T�6�p��b�#�y|�EHHXO������+<�0.Q��8~��-�%<ׇs]��XyB6��NVs�P�87��x*#�����a��EݍPT�O72�|~�s�Wm�];����m���ڡjĠTjp�1,n��_9V�?]��>[6�b�����"[E1.�r�
�����oD���V��[$i�0L�c7���'�A�q����35ɉtW$��R���0c���g�������e���U �N�ί��$�p��cbw�-�t6� ��sUҙ�l=�c+\N�SK�%7̰T� ��N�S`z��� �\�e�SfOT�3r���3c��R�2�J��u�啳��X���a�*��h�oh�[�3"F�6БcF
a5��&b2_I�0N�s�;%�����vB� 

/��[{-��[���}2Y��s���yP;*w�}{�����W[G	 ǡ�U����=(��i��_s������E��?�(\\�S��De�&~��ffMQ�D��x[Rcv���B ��%�(O��� G�M$6j���	��	,49f:�kg�/��f�&(h�``۹�~e���V#<���iŴ�}G�PIt��[����0��l�D�k�\Y��X}��~SA���������$Bf	�
ÿ��\H̾��ih�64�6eه��δ���w�*e�8�y(����&9��yx�B�"3y���Tg>shJ})h:���;s��/�r�տ����q��	'���  ��8,Q����A8�F��z�ON�C��c�%��b�'0륒v������s�}��� ��)$[�&��<�r��5B����U݂ڍ68e�?v"��j]׌$�8 ��q����-7���3�J�UL��h��Ю����G��.�� ΣR��a�}�V%KĽ�ȄEY���2R�\���)L��]����� �H����F��r����`��C�.Ag&R�K�F���8	��Ϋ���F	{B�Uy)[0����7)A?w�_�6��eI�;���4ݝ^h��>Q"��n;"�_.��_��":t�C�=��R��[���3Qp�X�`����c�d��u��,��_+3��d�|��E����_��О�+s�d�l����!ʈ)I����2 !�)���L�PrP~�� ��
Jc[��EԬE�{�A����&������;�ؘ)"k��e�h�L�,璱����_��Q��,r�%#�
�J
�X2�m?!T�;U|�/��L��26�h�a~A�̹
p��f��[f9��|��Z��e0A����$���-|B�����~�:��Dw��ГZ�7�N:�� $�蟜�����Xٽ�|�
,X!(���2�D  (��*	�+	��O����ti1vQ�p����z�:k����gFZ�ª�{�ހ��������=54&L�`�b���!#4iȭ̖ď���1�����p[{cFd��m��X�%;���m9F����Ӯx�����\2�DxH`@r(P%�EOY ׵-��M��[�/Nu��
Ӏ@���܈��e��BR�Z���r̭�b^���d���̟����k��v�F
���2��c�l�
���XoB�_À��e"^kɥ�#�*dǝ>����+2w�3��=z@%:~ [�6h`>�����(��~K�g^�q�-i +�&	$�q d��y,`[7P��o�z�����>��&�N��bx�. T�v:i����� ����G��$�M{xq��~���(wW���ɃǪ�~w��& ($1�A�w*p��wZ�����ʫ��,��PfxT�Ȫ�@n<�����rH�jKe�u�y�����Ƽ��q�������0@�B9r��@g�aR9=�L;'	>�2T�[��0�r�� 7��
Zw�cH54-��+@g�]?�,`��D�
\�1Cn�$�̬�".ⷖ�R�X�'fB~�n��"{�RD0�e��(oD4���N\Ջ�>�c��_֩� d��	A�C^*���`I��c����g�	��Z p^�c���K0�E �o����pJk��R�ޕvZWe�q��+��_�����/��
M;L},>k��g�_�v0*L����}Q�.���=�Y���-6�o�"�ȃ]W��Z+��J�ƹ}��
8����h��m��0�����
����ʔ��sqwĞ�cS[p{�*�N�v��ݖ�H0�ۜA��,Xr���D�x�c�Nm��U�T�������������82�L�愞� �1��$�7W�8MY�޻�u�2N�F�q������k�^t�O��0I��a��g0�_�"� ��ë�Aq$�8�
��2Y��d����:-F�f�ƨ�"��6����3w>�,����G�A�5�h�u��򙧗�1��"6<\CG��D�@DW
��;L$aap�"���5D��@>=(�-Y���	�PX���a�ým�E�U1�,�'+(tF�5���h�p�����|$��,��qw���q�gP4���y�(64$0`�Ʊ�ɾ!k�j�3�e&����n��7|�����ƈ[	��}�1��%�&�A�	���~h,���%�d@g,+L�xy}6R"AOw-����|2����!Me�X�ř�Q�& 3��CKM*�&��)�2�CQ�;0���/uҼ�\~W����p
C���f?�At���O�n�Z�/�\9{wQ�������}�{����P��2VR���0v���t�Rb֯����5'ݟ]tӜ8�;E=���oM�?�-)tL�x�Z쀡��� XL�X���|`��BG0F�xC�����������N_2n]���{*�`&�k3�5A/5>_�l��To����o�p�tr���3�� (�^uE0�	d6���ߟC�����h�6\<���:���#�� @3ff4{������@��
�Ã���_omt��n��`��4_�Ɣ4ma�ŜHX�P��hLf.�A�p��f���a���Nڿl͹H//��_κ_m���e�n��_��.���ⸯ���y��L��r&����(%j�U�w�R�BY"��?���O#w��,T�CJɒ�#(ؑ@�N8C~5xlR�0H�w���$����m&������ ��E�G[q� `]�I�H��6.=пĲ7�����y����)��7�e�B�c�B�m�w<y�ڕ�@x}|\�;���t�W�Ǩ���.�r��E�`���g�����rW�����"'Y��h�"8�� +��F�Y�dys��b���*�I/Y喆��i]�K�짖Pe�$��0E�Q��u�u���h��u�<I�G���e��BBB@�`ѡ�;|�<ٟ�qү_LE\�o��f���G�8�'/��D8U�%�M��ؖR����6��z�'	��޵8@<
��D�p.�/����v
7z��X�-Ǩ%+Ї��%rw|��ĩ
"0�*���f�ʃ��Fy0�ZO��:�VW�+��X��]�����ESb���8�����o�C��!Ih@Z&5���()�2H���$2� ;&���`��D��Rq�:\�Q��?c����L�+��7p��_H��(�!��AW)r��!>!��w;S��#��7܆S3Ⱥ������m���}/�x���:��-x�QFr�#���vd�?��G;�jv��{ֳ!���,K���^6��R�(@���pNи>N4'�;9���4,
r��x`�{ ;k�@�����V�6ߖ����D���vB2��I*B톀@_ĭ��î[����ӿ�3t�<�Z0��� ��!���ƒˬ�Ϗ�KN���J+9w"`�.ψ�ϊH������r�YA �5(h�A�i�!�m#�Mm�}N$�`\;�H�6<�ce>���/�bHE�6�M�WՓ�0	�8��|v"��`26,,<�D�e$�����RS�#t@��D��a4l��}��P�ȞN��
b�1��9@�G�I�!\J$ o�\Y��`�{��O,V�V����H����3e4���v�����;o�F��#��vœ���,��J� M�;-6[a��r��]�nM��F�P�{���=g�ѣ���ѱ�s_��V/I�G����?�ϝ�G��#&��V�';l=�o�kd+���Zѵ/�ȯ+o�G��M�B�nQb�k/�d9F	Ľ���㏣"Q ?����w�%�Z�Z1�89��@�cK�j@X��YZ/�"~ؑ9�<>�睚D�&㘷� ,e�<�>�ؑf��Ӣ��w�>�O���ުdOR�M���Ҿ[��/{yQU�=>_��L8m#@��{Ge�ftf�H���g)�flcN�9!m����M��
v��_�=M�v}�0�a�*̱��쬚֭_*�:������5�������HP/#�1�&c��~J1��#���	=қ��"���p0��iM��ؾk/������^]��A��]���F �m��)��V��:+�|7������Go�,p*6F�|�'��ļa����A&(�{�:�f,q��5���r1
>�ǂ���f굞���	�A�G\���f��^�\qI�C/< �h�����Ux���)�*���
Ʀ8<F%Sw�o����H�����(UԐikU�C��Z�gJʠXF��Iyr�V�,s���r�@ Ա��.��`2�8e_�9vi�+M	���Y��Y�Q':�����/����u��c�bڎȵ��$gp�oP�WжVղk�LA�C�H&-ob�5�No<�ܦ6N��n�1L�4������B���H�슩�o\��8����%��ѝAYY�l"�e��/�=���=aB�ȻT��G6�Ɲ|7�P�w�~Ɛ�Q�*K�c]eJj�%������r�1���{8[����	a"��SB���Εd�C�g&/�e��������!`��Q��+�_�n?I�|a����v��|Y��(�o	x��0��^���e�輖�����Ec`�X���z�7�v���f��n��$���v4J:�WJ4�J�H�\<�b����W�a��1�v��r�K
B�J�M9�\��}�6��P��b~�tB����� }	�e���l<�ߣ�r�c���||��f�`w�-�!���3"D$VcD0"ř+�K`���X-P?F��|8�Lt��)�6�/{}���v�V(����*��p)��D�O��`��en�P�GvN�"��u$4=��֊�vq�/�M����	3J���ڙ܊�*oo�r�P����:M|@��s���$�q���j��mUB���A��e�d*a��U�Qr�2�R1��,eN�i��L����]�ؔ�}�X��I�NS�pb��9#�:���B:"�k���W/�r_��C�^ׂ�t�-���m�?�$��3�lf �Q&�_Gn�{b�^_zh�'S��O�E�H�سׇ�|�s�a#~ ��0պ� W�Tf�3�I^��6q�����0���̓��i���(I���z@V�Z�(?��g�Q/{��q�tHA���$�3�ΐ�9��� |=�C�4e�N)��n�-��N���Go�
��&�x�Z�kJ=*jU<Q�Lu��s�����~�}֐�����z�6�~_A��I`!�u���:���^7�:ɡ�*_�
�q.
�`��%-����ق����H���\�����I�DC�oN9H� ��8���.�z5��/���!$	�;�X�k9��[�*�Յ��08-5u�/O����H1�s��_��б�*���#g}9�7�(���Ƙg��ѝ������t'��>��W	���67$�_$�
wX6���g��d�[ipwA�ܲK���(��_K�����_��(*[7IpD�����!I�w�c�p1wx%��M�����a��-�VYl���c޽" h.��zb����D���4Sq)��?�����з�l��,�D6S�+w�T�{m���b�S�ٖ�Jt��s������ԑ=�a.�w�@�H;M�`��pc�_ѽR^�"�� f���dZX���	 c�on�����CwDQլf�XIc�2����cQ�ɱ(F޵�7[��m6���M8F`�^r����a�jnZs��t�H*�$���C�@�0_�)�Cn���_l�!b�� ��Z���y��Hpތ��ڤ���%1/�!AQF(�wL`>&S0䃯�r�ѬH@,6!�F����qъ���+/��<YLX ԽW�̅x���_k"?谀�B���1G��������[ڝ*��VHy�D�~t$�*�L��rJM�h�̢�GIY��ie�, � 0X���Z]1��e xG��SQ���	kI,�&�64i� ､�=��m���=��d�	xq�iV���"�6P�Q�?���b�+m}�̾�	�w�w��f�� �J
V)��H$	X��w��
�$i'/52��BDN��G�
_~K��+[=�Wg;hH��!�t*�~W��1d\0�%@�sNV�(Z���VJB��B���;G���p>����+�(���Gς�������2��O��P��E��Ě��k����Û7�uc�/�8�b�ZWr��_&�6���������u�ʇ�E�j�Ğ	�L~�ب��&��j���Dʸ�ʹ��X&cʈ�JWF��;�>��4�z��;��:j�����>��`lW�d����&�M�v%!������h�B��_e)�$�n��x
�9(N8X-G���H b~W�U������0�V#�V޶�����)�-h�G�p;��3�Z�o��Mc�ן���w����<`��_��0b�
a�%h���S_�1y��	���V8���z���;���r�� 	�0*�ʣ�#�>�8�QSƣ��ఱ/(V3H��%IFzJJE9?��b�$w!��sd��&�aڨ/F��86�F^�描2�-z�f T��P(�V9����gI��<y�Qa<.�~[�N�- �3tƮI��<RQ�JMT{�t�>�Aޯ[�݂���D����萇;��J��H��G���ԛ�sD@�β��r�u�"�#�y�N��2�̠*��Mg6��(�b��.��?*jkK/D&�ޭLɒE��
�\�)L� �7�ח����loce��r�Ϡ��oO�L�*�0�N���Sd9�B�4�n_0i-A,���旧�e5�=8>u�)���Xv7n~��%��)�����gM��30��}����iL#�8!�r�� �)�ÿ��u���j��@�64C�%-n�?B� �Q�K�GA���
���5�9Xm�wAx��r�z<]�-��/��r�sP�$�مz�e���
����41��)�Wqv�/��"{lK�/��})��a�߹c4f�p���� �.�իzU���ZH�(O/����[y�]Հ��Z��:���������5���F)��\0g��(��	0&-�$H6w7�ѥ���Ԑ�D�h��b������	9��Z؁_u��$��F���o��\�̈́��QG�kϼ�b�x����X���0X���
�2y�n�&`ٍvu������G��{���Q����'D���[y���V�HD,�����S#�P���Eb�3wSm�����:��V��նVO���J��HmKK��FM�^�E][�-�2&��H����i��N�3R^PJ�~�5�ɗ�������f&����k!��N3,9�f�	1)2_����R���);�*H���U��%4&bw�՛��מ�������͑Q;o�j��h�� ������++Wl���^,����y3�}L)�BAX�X]B�pCiZX���h��r��v�����
��AE
��F@3E:������h����m�K�Ƿ# $	I���Ӗ��?�ޝz&�q�����Eq�?�ql�C<M�����`��ڂ���­��aOn�;��Ild�H�E�@%��g�a�!���G���}-���d�'���fP���HF���!&͓ZL�g& q$G �9} �Q�� �6���r��(�<��]Y�0�s�!}�t�<�
/�Bd�ʃ��P'j�ן���7�i?<\D#b���g�	Pa��Am�e�#��$!�O������~����D���o9�秂���W �P��E�	����%�t�L���S�W^_�怳�VHt���^@y� ��v����?�!G�C?}5'j�fg+��x����w�,z�ϜO-:C6<`@�B�a@(�kx����&3�����	a������[^jW[��v��ٌ��̍��td8q۹�H��%�������/���Ԥu&����|��$8� �k��4��+Hp�[��h[t*��
��Z�g�$�X��^'�3�7�lh�n�����-2f�����L.i �qo<�f�m��Ŧ�j���t�<����_/�ʂ2X�o�oPeJ�bn���RS��� �ėlq�]��������y}<��Ԗ�$�O���5�73B��)ڪ)�����58�% ��9��,85�п��HV_���g��[�ر�+�Q�(Wݰ��R�a�D
GuƎ!�o�'-����.�B��	��-��XU�`����@D�r��4����&��:(����t'��1�WL��a.�6��(��7ry���-&�CT���Rx�)uo�䍨��X�9}��Q@�7L��S;z��X��؆'�Wg�&=���P�AOCC\��a4�x�������W��+Qj�U����H~+�_�L�v�6�|N?���[�������,��s�����}T�W���8������HV(_�ތ<�+�S��b"��q�^���B8�k��k�E=݆���/�ģB�Cf3���B �^F[�@�u�W[:�f2��͠�_fnY��@���(�1�.���
��ۏ� �I/�P"���a�Yr���C笟�Z����
�@��C�*G�T�L+��W�[J)/��3��8Ys�[��wT�)k��������+�APk�b��v�o��U�F��2%��4T��}�ZNYk��l.am���OY?���k��aQA~
� "I�������9�?����hњ�a�a���MEI�.)w.�O�}�LoL��^���)6�4y�m\�˸!}&h�ğ>��1 v�,��mV���b��&u{t�^`�:_
����޽Vu�آ���O����/��G H�sؕ���/��K��/�_�r�������(������̾4���,gˡ��r�D��i��8Nu��l
l0��@v_>�U����Ta[U�� ?l����/w-V
�e�Y�7���O��&��-���eJUi�/��8p@��c��QWY$��`�|�,OB�������`�A)�'�z�A1:|�8�����_�u4��Y_e��|p��������#�t,@xW�[��@[�m�-e���/��TN?���f.4i�F�?�Ό$Sb���Z��&2Vŕ*	J��9�}��b�B�K�����atnуA0l	Ă%n�Xu:�d��4N����鰀# �u��hf�χ�zDk}��z<�A��"�/�zr����܁��1�B ��NlA�aMR%�<���IT��2�}����t�Y �evT����I��)� ����������=�X�c.Q��/%�@�J�Ö�9�Vܚ�3`%C ��<�}�`��]��5�F��-�Λ�ld�fJLi���wN��Eo�p�K�q�ɳ�s�Hݡ���e��ok}_��4�_s/�����q�/�-��_��+xq���-u)=��U��G�Wۼ���(���XaYl���q������l���`LI�H"0x�Z�1V��ey-s/�"z@8�����W��
��"�b��r��5䜔�:��5F��{���t߾����w�xCw�7.�,�)�m�o���0�T��`X`�l��(�ppW:� �^A���	4�Ԛ�k?���L�'O���$�c��}պ
�,2��܃�f}�`�B%��)���� >:a/�2B!�F/���>dD����<��`#���8ٍ���j���ܓ���[JH1��!ha���hq?S
t�c����`�$��?�d<4åW�?w����r����ߕ��1��g*�S�����~�&�lh�HG���?�Ql5sO���e�Ee�v:kSk�U���5��A��l�pye�z�d�������DG�kC98
_hKT��<e��y~뭢6������ 0t���P`Uz/F˶?>�g$pW�:K�ZEN���	`݊V_�V}��Fѩ/��9��z���H��i@& _f%���uU���!��q����)�
�}��qB��J�M�0es�Y+9-��.݆v{�U�E�60��U�J�b���_/������ 1[_�	�O�7��	��\����0P�X��c��z�&�o/&�on1�����.&ѯ��x��+v�<ۗ"6���� a<�|V�ǟ�K�&��m�`A(לA��p���ȒâF��!�+nX�<�X?���qږ�E���$k���8�����f�2�����Cg�*=h��NVb&����b�6V+f-��EM��6X"d>�Wq�����+A�����'��"}��/W�~�-����߽si;v]����_9U��V�x�Ec���(��ZJ<X��"���떭�S��ۋ�Ğ7�Mo�d�d�\X��y`�w�/�!�bJ5 ����433	�f�.p�8�bym��[�D��?ǹ�������1"ywx��F��u@���4D� �)�:�Ȣ��]����XJ�q-�,}S��"R��x@l�^k��4 ~=8���0�U�}�п̶�n�m�8G� D�n�*i��<��j�,��+䕯�q�jBi�҂_��o���b�w��\�S�I�4�t��f�_0�LR� �k���K�EI������m�P���d<<��H"�isq����I��񺠔>�z�CT��W���Ğ���؇_/�@�\�;�����YCe<�n��Ks���y����c��d��Gy~��Vq��n铔e�E�!Hf PٻX��x��q,aR��ry�1��@h��gt'Cm���ܴ�?���	�R�㲱�s�_�����ؼ�|;pK�v�~��+L���-�	E�v�ڄ�^w����
u5Bl���*E1�i�7��g��@^S��.�t���1�y�ȝ&�~_;��ÎB�2�9EE�(7ʁ)��ai�D(!c�a���ym���K��(���<` 6Ѹ�kO���]��@'�-k�v�
E�XZD*}��1���(�Z�������qL�%8(����y�ܠ�c�"�G_�[njFGOԹJ}�'Kܥn��>W� ;��9
_z�v��K�Dea1�p��Oev$I�N¶i4�d�H?�]��(��~iL�h�f"L{~�͕4���� �}S�a/��~_ol��%�3)q=�r{D)�aM�)̼�W��c3�K`*�e���e�
c:�Y��}򕴃�4f�_��k�kGC��ն/�����>��!R����2D_�bgH�\O2�	����ͥ8g$:#���Ӆ[�5�g��w���G�zF<<S3'UT@��/�gΑ�}쾩�B6�6�<N�b76��A6�����n��2�64H��J��gܾ���B�c�8q5��o�X�Ϗ��s�x#s�J��A9X����l;�o�.a@,ή��wF��n�a�0uTx��H���?��i��h�|���2�e$�֠u%�!󌕯�3[��6�ۜ�� ��~�t���4 l@�P}������G&���e�Qr�q�R�Q$�fI&�r�s�����"��}0��G	�Z�yD,go/�
d@���6*��͓����@�/�J!��!T�~Dֈ�bo��/�c�T�P(����lܝ��� �`�Κ;qi��c��=���Mf�p�[�o-�yQ\Qw}'O޽A���1�h���`�H2� ��OE(!\M�=�
)X��ȯLX�\�a��Q��`�a�s��5l<�f9GV��>�|�oʢ���	v��14��_e������`��.,�������\��;<�	߷�접&������Fs�$K;��h�������io)HfN�{�ȋN���n�Љe���M�3��[Ac����_C�]4��L��5̎�_�dY��hi$�;J��C��i�\Hiklp����Y-f��Z�F��ʳ�j����+����!�+}�è��.e��2�_����%�Ti/P�F��Rt�;>W����E���r���Ř�,�鎸-�����Y�f#A�}�k�� �u��.7�w�D�y���� ��?�WaWL~:L]E��U�>���̫���4�K�HB�zH?ƌ16������	O��F�0ഈ��u����`SS�3�J��L1�%�S����4/��q��-i����
�:���d�S�aA�Y~S��	h��vM�Wi�̕y���E5ջ?�2� ��6a�Y�MX�=�3Ŋ���j�Mc0�z�b�%*��L}}�/w�,�>_�齶����-�É
X\r�j	�T%��"Ŝ嵷[���_(I�d��1Ɗf�2��mp�U1�beRu�����;�b0r����'�B����m�bT�h�4�s>�h$(#�>��@��[����_M�E���+�W�F�,�.|_;��8%E�ʭQh�H�~?�	JοOh,,���"B��
�L�w����9���� �~qrN9h�=���4����FoG=+�H|6PslH>����vb����_�w��/f.�ݳnj_�q�p��Z�v�hJvhw۴�%I�5��Q��Q󐢶gԾ�cL (��i�$�L�֍���n�4�1�=��������v1x��0>fV.�a��DB�3��pN4�T���l�c�9<i�R^�ײ�e���Sv��)�i�W�&!��p�[���V�:��脗�D#�dp��v�����c���THO�N��~h���OE� e1ڌ銻�5���W��Ww~ ��'l|4�ЉYk��l�;�����L//�!B��Sx\���0F���#d�(�^g��J��x/rS���&�=�} ��@w��}�(�ɑw�Z��R�a5J��b-3��(7��_�^W�@���$���R�-r��B+�%�c�{L�mv�4���]�r���mK����E�JTr��a.��?�m��-L� ����r�țϽ�}��pȉު�0�,D�e� ŢĴ�z�j%^H��'�軕f}��\�$ӵ�Q�)��iǉ9w!�7�2���B/��Q)���yhj"��+eڶș��b�L3]#�EYY��~��hÃ�k�P?¢1��=tl?��I/��b��sP���7A1�D#"+�_M��tc#
����`Q9/�ɦ�>��pΑ䬦� ��9_C��͇ʹr�m�9�_�Z�|J���sO_<7�
;�% �[{@՗��'4_LU��&�E�d�{�,�/y}7۔^�
B�pۣ�T�Y��@���Z樱�38����b�݄�a bX�W80��J?wH�bf��}�`T���<'�=�t>�
�������/�	����#o�.�Fr8p1�d�Zn2-�0q��I1!���I_��@@�	�#�Vs��c�!Cv�o�]u�|��e�o�<K1%�w�Z���5�:D�|�ʐQ������KZ���d%���c��a�4�%�i�l/��.�)�D�a��Y�^���|g/��*��Qh�Ͽ{n��t�����M(��I�ُ��쭂Qu1��1���ҭWDK�"Nɂ>�m�lYXߺ��)��������h��o�G�=�^?�)��tk&ǺJ.V���(�-���l��h7����&�*�
a�_�pj��Pv>�F�Zg�[��}f��, �����Qf��'f��f)����,�!H$A���/�4���v���{��4�ٙ���N����2��N	3k���S��:��cFM���/ۧ�0�+1#��"6S�i�ׯό��
��oY��i������
��$��H�nHK/��0h-������D)���i� �;�x䏔�
��.۞n�_a`�����A�#���0���H�K$�U�هA �`*��_�T�e���Ϝ���	)��3���mh������#B��g�x�Q��±:^G�Lb���L�<%[�������6n5I�e�Ǟ��%E�i�`��H�**�2��D�Ĥ,$E1Z<f�����5X̭�s#�dۻ��Eg�gl	N��CcW����EE�����v����P�nb&�a�D��8y}�'�B4X�y9�	[��v�͎Ձ��=�I����D|���!��@��a*:��pD$�24zu�M� 6T�E��ǰ����2|�B��Tԗ�����m�6h�Q�\�߈ ��	K�����W:��S�Pɀ�>�����SC��dA5�!.o�_GԈ@6��}�ɗ��]���_ş2D:J7wL��e-tV=1#���l�)'���^�辊$GОӔ���!b�Ν�<�������1�p�ǻ��Ӌ�M��ce���%�����	�2�p�Lc;�ˏn~���&݊1��Q0���B���{��X���yN<z�_�,jn{m�����dA�Yq�V{��^�;k@�>�_ac���HHDZ꡺��������J��ǘ<��@�A�P*�] K�?/�eDtEoq�ƩT�� T,WN!d�e�O�=�\!�g�5I%��Ց���D�tƀ>H��Җ���=+oO��!�m�7+w��ӝ}y^�hF��<��鍘�q&]�D��8�"?U�����|����QP���}̿+��;�!mw���n�Gs�=��5[M�w����9�"�̦-{��)s(��B��P$}��,�O8�J�l��Om��:TM��C@��z+�m'��b=l�q��f���e������`;-�Nw�'������>�[�I�z�[9�;��퓐�"��[�?+�% �ە��m�M���oY��D�8C����[�J�9}g ��7Pb$�q/�L���S�ZH:��8�t!|�,	����nD�pǰ�6~e5���H3�9QJRy��bB��=F_ܽ� ��;�o'�A�%��/���`��g"��%�D���DW8��S�
8�삱�9��=�%��=��������w4�T�����T��9|�8q_q[���[�
Mِ�D8��
���m�<"<&��{��ZCz/�tF�p�V]��VܵJ�>��(Ƌٵ������x�b�׍zS�R��7�m���r�RY}��P��� �U�6݆�\&���͏�S���~��_�ڗ/�ӑ�3D���[)�
M��n��-}�U4?��o+��\Q��ܘ�ᢥf%�R��w���OdQ�Eh�|���-���JI�ۢ��*+춁�l%�T�k���َ4�|H��$P����c+2ov$�n�6��t�M��bѥ*\8�d[%i�g���=�)f��t����8�_r��}����婲��=1���'��"����]���ǘ��:2�KM�k���.��k��l�_�
��0�F|a�x�5ڊ�K�Ӆ�
)�齯�IŬd��M�����+b��6I������	:B
�ȗ"����0B�׆�*I����"l�o�'�
 ՝��c�tگ{���d�0H�$W��o���l�����o0��R��'�����JHe$j��4�-=���$_������]�ksp�*��\.52�MY�NS��'�o��=��~ُnwm��fۑ���e�.�'4�&H��	t��L���{��C���qY"v�}��K�S�hz�ŉ[��m'��XI�mńJ[�A�����6�)�ɺ		25��߂2\}�g,�%}|�W��̭L�ÆO�~�&���@�(��C�	�#�7�)����ĻմmSM6�{'m>�C���p:{��y	����tݡL�V����t��pv�}ąH Ad����&O�P�O�r�@TK�´����!�H�SI��(�!,�e�-7�f �%Z,��1�Ew}J��_Dd�$�w�J	��1Z:E��E�T�m):���r��v����E�*I�x�[d}��Ȥs_}���������L�}����6�63��=��<��������w�3�
��ŕ�y�v2�e�쬅B$�~�C��?ݘ��?bBE�]�v����ڿ���w2�e�� ����%6�v+@^_y�:��Z���3o�,��������H#Myy���rph�m|�X���a�o��en�h�wEK'"��U�^�ݡ����gg4���G��P����(.=W��v�W�>�t���<�Y�th������$	�3_�I��[��!���<��~?�B���*D5�CV�+�ފ��/�r� ����?s�
^��%~Z:��"~˗�[��J����%h�'�m�b><��k�y_+�y�H9#��3`�埐���sr�T��Gُ�����zo�Q����W��i����o���l�����"�S+�y-��O��ݔ�+݂��i�5x�i�"�)�$��͟����!lu�%9�l}�qt�����ig|���(�j3��]�ug�{��i:YYq�g��Zݶll3?؍��e/�[��d�M�����?;2��=lX�a��j��o��b]�yc���F��	?��m�tHĺ�pZWbEwV6;B��D��o��;���vu�C��B_9���ѽ��b�'�$����B�Q�'h ���f��D!���/��]m����e��F�D�l�������;(E�DHi���@r�ڹIi�ϼ${����͟���W��	�n����~e���$��]�'/���#m7��#����Q�������ّ�������/���w�9!4_z�o�����}9H5��Ĝ���GȤJgQ��Y}���L�=���yR~W߾_����dS��BW�����/�ZO��AԬ�n|ST�zγ��B ����X%"���R���]z�������}�)r���MP!x�V�}�F��Y�@>�~PBk��svv�+��I�Ο��A������}���𖂙���_�8�W��[�C��3}�tpߐA�ӗ���w;4	T����Y|Z�M�g���90"(0iec��Gg4t����TR�s�*�*+'B�����)�k߫�wH�i���'$�ޟ�� ���x��$���w%���Ǖ=�F/�&�	�31�;�Gۻ��L��*��}����*Ɔ/�]�s7�%�P4�����^��ʖI{J���l�e^<e�Ɍ�ʊI_/�*I7A_�߻8���c��^�.ZX�I�H�Z�D���@�������X<��Ae�n�����U�b2tT�(���v�9�3f�=r����r	�c2��ԫ�ڷ!ug'hP�Jg��e�{m�A:�N�JP�Y�����	�A����_m�[���-=��搇%�S�~k�L�ʛ�YskPJ���+��<h]�O~	.ƛ�m�Ӧ\&{����I�x�H� ;۠6�r>U�7/a���NR4ۢ�e�.\�)c���;�h��	��_wm�ؔRT�[Tߗܬ�2�-~M���I�1���e𛯙烫�A.�vI3U}�y}���V�l�_oj���0s�� q�Ik+���	�:1�m��y}&^�F)�|�N�W��D����8���nf-�ӥ[�&	7v& �&��-=f�h���ى����|�.R�0�eM�te��PN¿��,9}���_);H���/G�����C����_1^��n�>7�q����l�)~[k�2+>��~���X6��!-˟&�vO1�9[`��.q�����׷lC*��ܦ��e���Wd���.Ve��N�ö%���Yj������L_+� ��w{�$���;�]�I�q��_w��Ĕ�צ��=�G-�n�&���؍��lH���{��a�nQ���~ىJ>m���]���t鴟��c�D�D	oK�Ju��k̱�/�sʟ��֭�6�s~�l5Px�5�ܟ�AEv,.�ĸ-Hlg:�%*�	�Rc��>�۶lQ'�����4��UaNg�8�Օ�3�Dl��C,"�LI���4��/OB��c�	��x͚�ko��bU��Wӭ9�_�O9E�7����#U2\�#���)��2��r�-�\	�H���ÕT��!yF	Ǜ/��*a��#�����1�̳�@����1h:�J�xa��c�����&����tl>N3
�1�V�)=)�����}�y�'��Ε��j_�x������������74r�}��b4�'�tC{������7퓙���˖���l{�=�U+��@$D%ƙy���lr�B2e�$X������cm�u��z���VE��J�CGN���F��e��  ��a� �,`�#�S_bL;��1�/��w��=��z	X�XT !�>��j�c��K�f"�g���5%m?C@�?�}�[��5���y���.#���<e�*m�i��ee"i�&Z˵�{��2ps��&=H��v��m]�v�K��~9U�9&8�)��0!��B��<M>��C��H��$�u[P�?�O�r,����	O/�̀�(��i���J#�~9(\����mb�9�t_��C�󙸃�k?���7�l�sqy�0g�3�r�X~�xZ�6$�6;/���O��ūK�6��t�Ð@i�/�e�υ�N�y|Gg�'��B/= �E���\��&:1�K��;���(�e�#7�u����IDrVZ:a;��[��ܕ0`RT�/�n��9E	�t��j��h(�	�aĩ�g~�1�!<�E��T�ɬ�T,��b-�䀘�P?�٪m����X=�e�����T�aM����_Y�9��`��rl
�&�=F\LN��c-X��e@kY�/�FUpz�jL��.r��P�\�op�����X)�ܤG�g�`���P!��Oo>�'ѭ���$=N�[:t�y��% �!��N��]ؽE�2������Ģ�h�?�-��k�blW��I���+k����9Pa%���7��*碅o�����\����(	��G]�G�_���>�B� �J���]z,)�@M��;rN��ľs�,xd yP,�	���>���"@��f�>;�3����NyS�Zמ���^4����0�������04�A{ֲE&!�2G��@�$SE	7��T�)-H9i'�|��V���༒�V;��q[�����|�����&Cܿ�^���)�=�!w֫�5�s.,����v����J�������h��'s�i�����j��-��n��_G���G��#n�E �y�::�J^wG;S����s��n�6���%�9�L�	����wG]|"���6��P�� ����@�Z�����x`��,�ز$4૮;1�nيFר��W}�i�3���VqX0���E@sTa�z@[�M?/�Q{ |uV�͓� ^~O���yR7666�y�QNt��4�62���5O���tTx�x�?�w�s���xx퉜3<QPh6��v�zl��>L�~����e���ӏ�%����6:D�����cY���b��(YRSq���W���sN��ge������K��0tN~�I�^��y�e�m�v�3��s�)�����!�ֽ7-�����NH�Ye8`2��	���en4#~pKk+�����L��8�Ź��Ry���s��Z�����\V��<_]�{��j;�Ɯ�t���kD�����!��F]DnF�,M��.U�ѯ/��H�r�4=��f�?��ò����b���X���c�j��/�%Z���KwtchS�l�o�i�(-&�	�x�[&�ūT��^�N�p���Ә��� �â8+րJ$d
�^�0&��X��-���Rh�%�=��g��L�O��aśa�P �i����㨹&��/R>C�+��e;
�������޿3����Gf8T@Z�i��h Fz�חĈ$ $:=~Q�\ag���:����U�R&<�!�E��f_L�p�Sh���5��ʹlI��/��FYL�Z߈�n�۴�]ދ�S���Bp����2��eNv����:��)��v�}���,�x�淚ݩ)��J!a�8<i���𖂖�{G��.��0z��m�-m���e���L>�T�����"�o\><�}��ld��h$�p������>F�p��� �pY2��
E�t0�A"K-�1����;uȚ���$��E�e�% �C�ӌ�¬-b��;X�](�ܧp���p~�S U��_	y1�zQ�\��{6�*5��}\�N2��ГpKe���f.�����	�/��?#���Œ{�H����t��.O��ns��q�Kb.���@郍(>�/�,Z���6���S�*�3(�&°�"�b���1[>.Fm= @*��-1�lf���bp�h�S�ڻT�!����P�H�M�;{+*���zc��	�̣�9�m�6�l|yk�jO"T�n������_v�fK7��s�>Ǚ/)���v���V�l''���6�eݻ��6��m�#����ϗ�$@J�gQ[��[�lk�j~�Rl 7�,������◡�$c��m�C���~����ܺfZ�R��-�hM�Z�~I�tE���BjbJJSAQ`(	7]��Mf�I>��4�+���=M	�-����w�c��ˀ�h��
��i�2
�Q����
��U�&w���ܩ�sQ�%�Yu�P�� <�ًDE�F��G��sޅ���C�� `P�:
6�+!XZ�HY���3��k�h(P�T*��i��Fy�Ɵ�!	����ݥ�( W6[T�Q/Gc��#��s��:��>���$� �Vح�i}��a/�� d�#����Cy"<}ߒ�Pǎ��A�^Z���-
RP�k��S�/%�f�Lt/=*�w�ZqCUڠ��L8�zL@�Y/�X�X&2Upw�D�#���om���Ŧ�	?6������Ї>z���	s�I;?�P��kG낰��h�Z^�Yo�!�����۵.%=�$J������a~��g�q�����e�x�6��{���6���Jd��C�#]��)�+
�e��qO8ؤ0���݈�qc\"U��|#�ݢ!|�qě*�t��d�M5�CH�������1h��&�vC����Ѧ�H��o]X�=�Y�U0�}�Y`���>_��b�['s�{��`G����e�B��]�抜Fw����c(�;:��=/�!aYN#�>��o�R��Y0�H���j��.^L��gh����kВ5�>��c�*�J�k me��h�?�UI�=��_��>�2=��#�У��P�\���3�j�B/9�/���>�pJ��O�e�ہ�kC\9(�p)1�Ta9�[�.oT��Վ����'��
-�S�]�������*Ǹ)��+�١�
̻���He�pe7���s3�:a��x��Oi�7DAwB��@�[����jO�!��ؽ$[b$��o�<E�
�bq��[��軄dd�a1�«��)}��8�d��׉(�a,
>,�:�i����Iˬ���/��qe(xJѢ�;\Pm��k8�C�iT!������*����>���EY�'�g��7���B�����^\6_ب��'����@R�P�ZzGG�.b_Iu �>�_1��i*$IV7�7}���7I"O_��%-�,渴Y�Ch�I�`���Jl�$4Yi��)?[�×Æ�.4,Q����d��OZ'�2��D%|�]�&���(XHM�~��|㋑����Ѷf��`�U����"W����42GI� `��6;^�=_���3�P;^]7����\��H&:Ieb%�eӯ"����x}j%�(@"�۱[��1���M�	�D
����B�!� �6�,.X���Dx��C��._�QTF>��
	(f+}_���?�;±�Ŕ�~n���*��CZ)V�a�+�_�H_c����UT����q}'��xK�q_/Ӊh�����O�FVwcm��k���1c�l�l�tf����_��N�g��7�C�Gۢ0�#ӗ������m'��I����B���G8��<"�`��+�땎
E�St��C`�8��A��V�(��s����K�}�ؑA�����!��N��<eWxw� �6����k���l�8%�^�f�?�}.�=D����1/!�'��W�y I�۱��	�E�ϱ��|��Qe�D����KIM��/������+���}�����fY��3�v=�f<*<* �>fI��h_�ӃZ?�|x���AB�p�!�[�����#�xF0�7�}���G�z��b4A��ƿ=٘�Pkd��GX���Jݒ�����_F�a6��g�)��#�b'4V0X �>aw.�6d��v�t��,��<'�#	��ۍz�#�5E�sY	k��	��1*Ef?]�SI����G�λץ~;q��:9�x�CB�X�Lz8FN�,+�E_̇�$u�_(�N!F[��9��Uu��>?��S�^�_��}S��_�������v�5b!A�����2o��6mٌB	�*�w���!�4���M�צ"B�\0����*4���\*6Ȍ�݀֝6P�o��!3��Dg@�EDLX�z�*��=|ZTGT��x��1�TVtS�`�U�%��f'��H�^��(Ɯ��a�M��!�:�*Dݴġ�/h`(��n�CAC���������A"��w��527�s�8���AC��wm����W/��h��Mf|�d�v����DV�B��k\@���Ƅ�=}h��s���<V+ޓ����cFEbN"�V�lC������Ã�D,�p�����ϕ�ݗ��7qZH���;f�wB��\4(_�DO�R����(�<Hҟ���N2�#����\SJJ�/�,��]�-�����zީ�_�����PF�ID�B;�a��ml����#�ϭa�ڂp!��)��7;l��
4w_����w/|{�{�9�^)�zO]:b3��M�٠��F%��܎��n 83���8�LqT�#�b��t>����TY�9P�x�D�=)�`�>��%�s��s������aZÆ��'t�l�/��ޏ+Ww��'�$MSh��=�3!�3��rWM;�Է�,3��(7X0�PL�Ō�@0A�3R@1u�$������s��N*_"������*~n�����/�3bE�����1��xƓ����\߇��%��K����X�a�[�#y�F���
��"'p@uye��k��@�L�2t%�����ц)�hA����ޛf�΅�o�؃��:�Y}��E�!�1/��l�K��G�6~ژHPI�I�6��F����R�;R���M��1Ԟ��g�/PNGp��Ea�~�w/��@�S�O��Ѣ���g��1�N!`'x}Y꾴�}�w���Oށ�gƨvCc��ҷ(�se."B�/�l�vò�a1�@_J~�zx���D�2vD)�d����YP�m$S]�,��mv,*q�����|2D�ϳ��J����0�E}�A����wuQ��� ����)�C�Z"�1��pv�,e	�|�Сӟjk�*/����F�1֩Qb
n�Xp*X${��Y�A�����V��^_www���hm�X��w�%/��T�Y�r���5S�4;8G�#N��I���Sc�T_ �c�l&Jb�_?!XTt���2�΄X���2ߔc���wf���s�	��ҾY}�i0䴦��ʝ"����/�ި�M6��$Cb	8`^�p@ʊ_�zn�)��룝y��Z)lI���8�I����ѝ���+�	��q�����יs�2bShr�jx߹L�-�_�E��זl �J�
4i'�Cd�B["��o��5��N%�_5ɰ��X�}ZM!��*�C�[MX�M,(UK���2���g��:��YB�8ǻ/c��ǠO��@��eHr���Dl�p/,O��n[�� \t�j� �d�/��dd��Иm��(��c�G�DQ��d%~0�e*c�P�G��D�`�[tU����{��;� ?��%|f��>��*˒��s�d��A#s�l72�ڭ��Ѵe���0����X���r}|�c��*�(��}��O/�%��$�J��ȥ��%^S�|�G��a�~f�ʁkV~g0���7,3��Z4�u�ZN�aS�r��@�j7GBL�� t&N�Y~����Ȕ�nbن���(,j��د�������p�4ν�h���a��9�7u���,9/c�=A��H����;�M�k ��aցh40����c�a���������H�g�����(��{�(��v~HW�����A���۶�G�բYiT�g��|�9o|�˹Xя�c(tD HZ������eˆľ$1��BL<�Z�����0�n4�:}+"zV��@�b�?ݻ��El�`�QX+	�u��mǄl�c��_l�FCl�t�XTM]�/V��ʨ��7��N$�s����BX���o���-;�˦��`�9q���&���	B.�=�t7�me�"��_1$f�	��E�I�ĕ˟��r��p\�MV�P�&<�,��/�НQX�X�ǉ��Ձ�`/�=�s�`z��h��T�Cr}4�Fvd��(7<|�}�ͩ-�m{�rb{�;����{L_/�eN1?��.1�v�M��+��$E�	��Y��&�S%�Ym�Qhoㄻ���e����I�Ԋ,�4����P��i%Ԉ����];g�E
�WS�ľ]t70��X�t����|ew���o4�W:��Ǡo3F��؈�p,�!
��w�
�:�׊[`�Mݎ�"����n�w7W;:���z@MR��ܘ�X��(� �����?*A�6A�3v_B��
".Aɹ9"�����%�%J�V�g�$��L���"���Y�VI
�1p�DU%�U̹!��O��ٙ�s���/��Dlp@$|����B�c�K�v2
]*�b�0���e</�y��R<��$-��.��"V��4�����o� �[g�k���/�^�ū�B���	|�J0��Y���r�נ��& 4(�>�
�$@�����'%���AF,X�aU�b����&\�~�]g$0{?4��$<B�A'�����ԙ�p@>�w=���>���%�����nA?���b���D`��[Ƣo��@���T~��G2HV�k�;hT�fӠ�{{&딋m�yE{���k���~o�#;�;��p��y��G� �C�s��O���+D1̾�+���5���O*�����nW���݄�C�U��+;�P�F�Of��տ���qKg%=жS�((R����Ý�J&WC���hZq�Gj�:�ޏ-��0�vG�f��E1�o�A������+˅�}{��8�%���ʅ[;���+	�_ hH` ��P��?��p��p=��c?��p\.����Eu1����hD���z�MJ=x���H�|%���u�������*�PC��:�ZD&�����WtK�hA a�ʇ��	��E��~எo�!��3I�S�H�9�����⧨a��wv�����hA��tI9����D�n>������옮���|�%	�8��u [KX�Q.$�G#�CX���/W�#��j���"
��"Kp�o�bi���;/��~��N�t�"���2E�[!�va���v�()(�a�lg,��"��~!�f�k2G�+5��0���!�1ܻc�Zj(J��}@�Ј�}�t�a�����.���j�3(�;�����]�ɏ���"RҺL�������6A 0Ge��O-�/̜=�0@h�Z%��M���N=Q��e�BG<��)??dح#�Rb_<H@�ݪ^	����B�w�|,87�aD��vǢ�/�`�����A�m�AG�kn��`�$Wv������_oվ�#zd�>�w��ÂO�?�h�?��D���q}h�Ap�VKT5s�M���A�/�]YH0>�� z.�U�]�.���2.k���j,(,�\Q��Z��sk�*KJ� ^���*�H^�z��*2vp��6�lk�-7�ۗ�1Y1�=������֝��}Q�A&��K�-���.vZe�jOyr�2,��o��TD v7wtWv��:,��d�{��eF�fO|�������x?��PLC����������K�{@q��.((�}�����?vE!���̚��>
u݈���߈T���4da��g�0w�(���;�!�2c�$FX��!�}�@�����Re�JCE�AX��Fd�,]�we���7h���5ۂ���T��04$����,��Pݲ�/������$x�ˉ5���R|X���+˃y��5�6�謞�_
���H����DF$&��	�S3��D��LPG=����{:$���&k�-y�8H_n����ߍ�w�J.�����>�� ǣ��/�&cJ(���-w6�0�Y �i�M5��7z�x�_�%����L=�#���-��hr�h�=����(7>[�l?�t��xT���]��8��ǖaQǯ殅�b�x�"̾�!���6�����Bw�۶�P{:Z:��]�����m������Ѱ��^��]Rwl?��'-lo�,��pV�
X}�l4��x������:nf֟��H���)��m�nv�픷DWF��
̨dF��@��J!SEP6A:�3e����|�F�yX����A7
���ϊ�L��ʨ��	�'ފ>
�eI�s݃��yj�M������w�P�e�b���t�����#r��V�=�UZHW[EN2�s�.��0�N$V��-����PNw�ù���^$�_!"�|�;+��$c<z��upD���/��2�a����_�.���F���정7!b��@���m�����ɻ�R/����i��W��2���������dU�ȁ���!���D�
�h�#�y���U1}��=��A���l�i?�&MT2�2��#@�.$�F�gXQ]�X�&1MI��S��d�-�^�+���m|����֓<�A��˗{2�r�V_Ք7������z_��?���ǖ69�$^
���H�U��/xC�f_M��Q�BG�W%°ֵ���E����qE:98��%1��/��c�`$no��aW\`��!��h�g��<�g4
�G�Sغ�]����	9vi����:��x�8��VFV���D/q�^j��'���f*�/��Dab�%?�����Th�TD�ZĎ�]�#9��G>׃$zO��ܺ��=���;)XP,��Y%z�g�SHl�P���u?Ai៿�Ǡ��'OC�q���<:0�a�EK��K�������Jƪ~ؽM'G|�{k�/oe.���L�k�A�.�~�ĄV�f��C���v��β���K.�c����_?id����G�l�{�$s�V�m�߆�o>Kދ���oe����"�2�5Ѣn}���f3����?�xJ�T-��.K�x$����`��FH�0�P��/�}�M��<[SQHw���=2=�E̾r	 I���3O�n�z�١ �`�M��i�a�$�o|5��r��I᾵���}��w4i���d�vq�_��Or��+/���qC	H&��<�jpa�S+� �t?)0�ý���.LT��N~h`!��o�� �T|��v�l�#���
k2�\B����[���&��?׾���&�$(�1Lh�l���9���N�`'�	�6���ȯM.`�K��R%�|H�j~[��ġIPP	 u�n޽z�NY��__5���aM�� {q���H� C;��S�D��J�0�� �sG0�`�1hcPZK�C/��gI{�J��	��m9�o���ݖJߍ�K�|����{�1ws�=e�r��\��W��e�%��g�m�'�ܙ�� $��r��
�qZ'���-�G��������,M��A�z"���/Ř`����>:���2%�{��[	|i�	 B�F����������rמUx΁sm�����x߷&bY��}��d�
�4���jnZ
�1�:�k"�P?�YiľC���������O��g)���A%�zN���n�ZW��1�W,@��w<ޑ�A*�!�<�~���`��'�Y�H8r���gċr�w>?/���Q����∕���	XǠ�X�{|6�7�� �1h��K����k�}�u~�/>9Kh���nЫ���x�h��ח��r���p������Q��f�rm�e�?��XpD�X�|E8�y��f���V�J�Dc7��H���t�����X��򘸭�w�Y�������i3|�ӹT���̩��&�	x$=[r�/��Ăg�����l�@V
�6�;�t�h�:������Ss�A�1���~w���5g�̤�8OSC��Mf����eb+k�����c���˷�C�e.���~�v_H$$-�n&%���}$N��줩,���?�L�F鿬>�9P�#�h�|\�l�P�:ZH���
&�Y�5N��^�x(�L�SڟpUR��8�bs�V]q��>��|HΎ�da�o��8җ����&	�jjc�[2��2ʅ���]�dlv���:�G�������~��^��l���*!�v�4�L��W5�>6�Q�u����+;��+ \u6��+�ʓ�-7�w�`���`���D�W��p��[#���R�������(�#Q�.�ܱ�m�
��il�������2(R	
ˊ���i+��&J�O�aqF�=�u2����F4H��B>�.�_P���c��Uc�`X�n�rt&�p���c��Ê��8P]��6C��5l�0���a"�jhg0�s��������2\�>����@�7[42�n�y�kѶ�_ZL�
X����k��ݿш8`�Aݧ���,�&%�f&5�tG�,r�����w2�*N��M�o���y ��X]�/�vP�m[���;ʑ~��{q^������#^���7�zK�:]R�+�[|`�����7��q~$td�튕��$��x�[��r���tp���ҫ&+HW�]=�N��5��Y������ �I��}1a �g�U�
��ĕ31�8�б���Sm�Ⲡ����h�A Lx�����l��d%e&w>�/7�O��_D ʡ��Ak-
"�� |y#q��s�n�lQ�⁺���+�d���(����#et?͜Nc��k���2��"A!.����~��Z�������b��zX�wM�}ڴ0&+��ٔ�/�"������;L��0�2V{4���e{�G�\5e6�;fa����A$x��GW|Y��k �Lb�$W�bcb�n�q��".R��[Avz��jJ���&�:1��;8؂��|�U���gL4!�^hX�_L�����-����"�;m��}�JZI�l�8�VO=���M��n��"�9Aq��C
(݁�p�Ua�����+m	�b��]
��0����0�P�2�>_8`�BS�3V�-t��i�m���P�g4S\x�"��ܾ0���b��n7��o/N���
�N:�>�%�,k��YX� *9v�{������(5(r|i�E��s�&P�9���c3�D��i�NtH�1z�g~��_C�AKb:D����{��f-i�=[m?�����0�`F���J��O`���i0��^�a��8�˘ٶ��_�|C������7�'���۶d�!q<��,.%�ױ����2��ÉҾ����f;�.>0~3�t̙~߰H�Yz�������������P�1,��Ks0����!��|�����^�Bl�{q._R�:l������5 �>_0�aD(�S�돂>��Z�ܟѻl<�(`�QF���`��r��!���5�"�#XR5��g�핎Wܣ-��'��9�A	Evq�(��1�g�JՎ!�V:f8m���+��t����et?���0��|�44?c\o����-����I�7�$$7� 	&c�%5�l4<h�W	�ɹ�b<���n�t�d��O���a�:@��a�&���	������Ֆ0��v�����|��y�ڬ��8��,F�A�����_�Bf3B)�b������fBb�s�FO�'T���Ai���ac���ږ�;�w��Dn��9�Nc�s���P��=l�W���2:.����>����eA��#�x���~[�%}	O�����G�s�<I3A���q�`F
<4�TD�6�`O���<v^�4�'zV�H!y�N���
=}+��W}��r�a��/�~�>$[�҇7f���\k:F���(��Ŕ4L�Er�)�YZ��
 ���_M?/�\�}�AJ1����9�/!�vP\L����8���l4�/�Կ���PS�\��cvI���षvϏϏX���B���s�%�̚Ύ���K �G��%�Vl�Ա�|o�Z��p���qm�'!���*�B�jm�ϟ���.�G���n��̾����Ү��윽n�y�������{�����O��=�"���9�	�<��,�)Ut�͖C���m���_:�o�/����5[/�K:!��c�cNvA�zKM��HܥRB���8�(!����#��؏â��c4.ͬ�	&�3ȸ�Ra0���=0m��Yn��e���Ɖ�=�Ȕ7�sa`F-�݁�ԓ�����=��Ax#�d����"�ɄJ��`��x� �w��Ċ.���}4ߜPl'���5�?`��H�l傁�gj�Y�=���_h��Vw9l~�%����t��A��x47Kp���e!'����ܣ��7��a������(��������c?n���������q��2���5 �&cYx�a�ԗ�0HM*F�m�j��HX�X|�Ίs$��ii�ӁMDxKm���2.t6�O��*5ծ�͍�C�dσN�9� �������D+�8l��}�r�������ln5&=�Crq�b�"`��/AY}��Shq\�}
�%�Ի&�m�`\<�k����v�y��$���+߹�-����u��c���E�f/������24Ғ�t�� 	k+E-I�@��M{�zq���8���yο�$~����Q�)B��䮏²�in��in5�ap��X��u~���|��b[O�|<��R��U� �����cuue�0�E ���E���p��}yt�ĵv_��RAv�H�"���wJsj��_&�u\���+�{E�C��վ�!,��"<����	��ޝ�%٤����9�Г%�a?�������~�������z�q��th%V�����/�_-���;�<Io,'��� ������1AКA�P�!`��"��R@�@'8�����l��C�Wp A�#ǣ�/�Oa� �x,�uSiˉmH{O���/����ͷ��v`\����:�%�hC8��i!�)�	�b٩A1q�פɩ��|@R4k!#I��3Zمp\
�G���5�~黹�_A��D�A8֖��l3�`���,��`�6��F���郪'�A�f�h�7v�E��ǴF� ia%���It/�Et�M�ڕ#կ�H���%&H�����X@�}o�w�%	K����Y��ش늜o��4Ȇ�H8��R~\��8��8U4�ګ��j�>gX�#��.��c}��s{��1Dp���#j�,)�:���Y�;f�Q硽�GeC]��P�ֆ����w�m��T���g�P�K�� �6/��#�	Z�q*t_���FQ��N�������@�~���ƿs��;y�6��q��'\�Ώ����0��%<�Z�'�}���/�bE46��h���r���d�X���X�͕�\���*n�����#(&�s��t�en��>��6�r��"�ɏ�a��?�V,�82h��������$Fz}�a6�ِ�@[a�	�F��c�㯷ORa;�?�g�����U��?=p�G?��N_:�<�l��(\v�Ft��Ƒ1E��s����ւu��~cY}��[����M�8�rA��inA���bC���V:��A~D���n%1 ���[ᑟY�����^���'sgo��,�X���3���Gv�pR ��v�����̂��X�� ��q]N+>Iɒ�%�F��.����Db�]M�~� ��X��
��^DA�	�nG����)�_����2�s�k���Qg ����ܲ'
�Q��{�R���AyDHC�A�ut%qO
�{�!�$��+-[fRY�xW�{
+���OtO-������r��"-cF]�V��/���H�rC8��<8�V����"��������&r�<��1F�y_�;�F����۶\ʙ}���pBy�����^aO+��||���Թ��ؑ��:v�Ie��Ge�ԡ�@�_������xA/ҿ`O���Aoo�LP��ײ���D,��V^a��!��)rC��@��7��M��rƾ]i�[#(Jݽc��ce���]R�xr9��D�!mdC���9�>	�[�<��<��w�*�4m�|yEt��D�F��C���(�6F2M�44wA/nL^3��T}ﰠ$�����+!@��,�\�������)V��a� �g$�毙��Z�iȵ�#�4���R�X���ǗK�w尣��.0 89|  �G�FÃ5]�G���\w���ΈV��Zc��-}��D���}���, 8xY���3�Kgr�d#m=l�,�%hڟ���i��%�>��O� �� ��Z��p@sܓr��}ў8�_9�e!AIh����͹�26^&�}��JLR�U�L;d[�ߔd�G�[&!�z�O�|��D�Dў��m��Wl�v�j�A)��#V�7��X�3��nk�ѡU�` �O��R?]�[(R]p;e<�W[���<{\��F���
��"|e�@}�<�E4���t�.j��q�����>%���HI�4e�,5�n�K&X���a+0h� ��/���\��.[��<}2o/��"��������g����wK�FIR7����[�)�m�^�>\K�Ȕ�+��ێ�r7�T���N��C��=RS�@ޞ�N�N��k����h:��`�-�w17����ܑ:	A@^�*d��%��q6}Ɗ?���{��P���2�Ǯ���n���3���
��	��lSu������>_��Պ�+���6T9q�o��դ�溽[����;�ш��{wl�X�#��`[v�A�5y'Y��J��K���s���n�m��9|6�Ñ�8���{#�Lw��m~_�v�6��p��+?���e��u�%�>Rwm��v�Ү.����<s��$�笟š��/��8�"L����V�i^����/�=�HP"0 H����|@w�� %�_�yOm��_�34���YRW�e�MAT���wX>3��Rf��AcAK(a��ן(��`&h���󲐣}��a9b�����c(��dr�}oK��,'bB��g/�����E�i�b8&�1#�äP�6l|��O4�Ʋ�|l����3�]2�=Z��u����yvw�Ծ:D8�(&�`g���L��iv~%��W~t�f]4#�
7	�����Dj��2&f7v�͹`�\~�M�A�bT
��1��~睭�Бa�Z<-K���T����)�b���dB��N8��2���FqA�g����$�0��3��j4��H��~^H�m^M�,�<��+*1mک���As���!�fu�n�8"��"d�/���2� $(D- ̖F�о*��;	]]v��C���*J=�q�t-?/�)� �.�?u�j����5|�ٓ\T��0���./xaJ6!o�0�Z:�ߏ��[��A8��f&S��jK	�K�e����44��)���ȯ��0��'n�B�����
S���Q�q���5$����l�� ��lC�g�W�Y_d�2õ@h����%\sx�ך�*�AU�Q��żE�U<�Zq��ːjPX���sw��f9J�	���})��k�FI	޲A��%���-�2�����׵�d��M�7�/��ۘ@��5����?�x�6:?�<�q�b[8���	fs�7���r%n0���K��	���z:g�|&*���J���)M?�4�u�߃�R��t��¤2�5N�]��{����+�� {9�����3yo�:���b�rp&7��G+�#���g��P%c֖�e��&�g��zڠ���}r�ĐH@,4y����]U7���w(�`�/�SѾ��"��! ����証rj�;�E%���/��-�(�C�HC�yR��_e>7(ٺ<t�pD(��s��Img��|^�
����!+4���}�w�B�Ю�S���=>_��v��<2�vS�]ޑ(�'9�j�q�Z�n�-Vq�{��Ȓ���F�����n�s.u�ؔ�����׾w}Ͽ���$Fu{�\^�,�=i�۴��e�{��q���r(�Q������U0}N�8=0
V�b����T�!�`����+����3��@��o��
��s�B� �Zao=6,m7K�Ww> Ci�='�j��0�1��b=�^�������o�7��T���\Ǳ>�1�	�Nۙ��������PU�^�O�
��2̥ �W���"b�0
:�o��hX!Q�*�Ϫ)���f��'�f�j����X:�G �&��,� -9�Υ��@�ӌ8.-�4'��wY|�Eʂw�n�Tq�^���޸��F*jS�(��߆��.�̾��\^>��2P��	���i�ۦ1
�K�o[�{�[R(:�h�_a&BጾS�$�
�;ܲc%����?)����Q�Ev+�{����G��o��0�D�J\m���yDr�u�������h�Rhq�l�~Փ����ǚ�s_�����N���2хB@U��V�������	9�;x7��)|&e�q�@-LN�4z�WM�p(�����S�c��ͩ�`�c-�4z� ִ��f�2�x�|r_�$i6��L�o��l���SM�=�����0S@�������L�͗m1��e��l� H�'!P��ƻ��lK\A�؄}O<*� ����X��hũϦ�M���C���0OE޾x��~��;a��h�
WpTe�4��/�۳�,�&:E-!�����"@�~�Aq�2�m6_���qH�b O��n��S����5t�'�u�1�3E�?M_�(")�]�t������FQh܎��	��NھAGł�"Il9#�si&� TKu;�Z%��-��
���$9]��L�C��	PB�ǹۉ5C�ڢe�%���ck[�\�8��@����8�D���R7�����<[#ē��SI={2˩m����V^Q�8��0F�C6�����C>X8�{��/,O[��������e�}˼��ewCײ�R��Pb�.&X9pQ�ŝ�D�����ľ����'��
Y���A��j'b�R�B���R���c���: ۇ�W�#N\J��A���|�|�n���Xi1[;�`*�pƃ��X���Dj���)8g/<�uB�Y(_T�!�j/��gq���L#	O��;�B����Q�Ћv���5��Hed��fAny��\c�'/�R �/��CJ�v5܍��U��B̊���]R�t��Oa ��+������2���`^��%)�\����w��t+�𨀘�q�I�
����+��v�j�wb8Ӎ��^G=|�T��[���=� ��o/�HQ#���ߗ3�?�(��cC>�s�;,@!ArB��
�>7�~_c��&PN9�[n�����
�B�[�ܠ�c&#|�X�����ѡT��6L�ߗċ2	
L`Xg�A�Zu�Vy�R�X=n#�=+��bP-��+��\_���tF0��H�i}++l
~ҥ����<� ��d7������h �wދ#�m�'�Z�F���������Q!��گ�WHs^x����<�,Jv�8�@���ѻBE�D����B掴%@��F �ܰ|�c��^���ԯ�k��o�,�s��ن}Yj:�q�L�����I[/�@�"r�"i%���hVꀟ�(�1l��Yz�m��j��Ќ��X9�O��&Uz�&i�p��jNDSz�*y㉛y��/��$��� �S������`��E�G�߇��iZ���nA��b�Y����'�A�p2DA�r��F��.�9e�w�/��b�L4��1��Һe���<����K�k��\-�ȇsw�
�3U��Xb�I�b_����J9|�L��Fly`���W����|�l�%]�ଙ�z��|"y0�3#uY��]b�?y�;���4���VaP�N���ř�>z���B/�p#���<�lϙ���/���8ݕ!��_R�.�/C�.�Ai9u(A�K�{6_-�$j�l��a�	�~軂��F��Ȱ�\#s�իc�G1�(��	������m�H��Bq�z��akCup�=օ��!ͽ�NʜW����I��_őh�,�/���Z�8����6�KcE�v�⻏�ɸh�&
���R̕�x����|�G��15b\��q� ��^J�����0y����I�{�w�<��p�� �R�wF�ࡰ�+r�!#��B�t~�]e���u���%�p1�J'���y!��Aes�l�0E�8�2K�du��/�a�ՅZ���;���
b�qF�Y�����&��p�X������t�!膎��� ����T���<-� �gdI4�qO��"�6�*dj�c�,:���A����Q �`�� ��Q �"�=2�u���)�뛇Q��t��X�����j�_��u��d[�ղ�8&�3u��+ZS��}�S8�ƅF��[���l�1��LN��o�q����%c�x���;�ɲ�wb�����/�N��n��nD-�:����i�r��e�X H(�E�}gS�a�믨KI����.L��z��~��h��e�����cܤr<�A$]�Nq���bV��i��S���|P�<4#��� ��9�}�r�ćl<$A�=�v��Pe�UWYZ,l� Tkr�)f@YF�������wX���OY~ �L��j�<�E��0�U�CS������!
	�P�I�;��Q���jm�؜:�W��� TP�rF�e�b�L���֙�e����'
Wһ��ۻa��yX6�N��u�;��qA!!���<��癵���;"�2��B�C�)�mnp�4��2o�j������r�����y�v_fCBf��I��`��D���m+��FJ�/�t��lQ�˹jc/A���n�ymJ�N�� ��Ѐ\),v�[�����3���(���Ƥ�~%��_1[i�� ���r��l'*�����BzX�S:
_��l��AA�3+	���q���A��7���6Nc�QP#GYe�/��n�C�*G[.g����q�9e�Hf�b��Oڡ����+0�J%��;L�/&� ��AaܓE�o��M���ǿ�6�|(:�DW%�p4e�pGY~B���T���@����E	��� ���)���=CL5Dh���x��uN���.�4﯂����۔`�ү�� {y�)�C����D�.='�7w)ٰ7�v�:w\b�{����]�t�����s�N�3m�w�� 	��V�X"��%N��**��I�t�/���k|5�}#��H[V,쿸0e��Iobt7	 T�7D���"��u��W~_r[�c��?�����H�7'h������H����nD��v�Y�⅜���O�w��J�NT�!M��d�8t'/�d64ʊ�5�I�f^0@�K0����f1�p�w#V>������/�6s�+�)�N��wq�ݎ����������~>%�P���O����oAАu��:H�	m��ήgE��{l83�m�@��0�ߗ��ABD�o�7�d 7�w���ʫX��ڢ�X��%2�&Kͩ�&������� !�@��L��3�N�څU��?TI�zS\q�6TA@����ԗm��h4���e�V.%AF�O�w�{�w�����]�-������Zp�D���ᖶΉ=��L�.c�:�bQo"��
���\E]�a�FJW�-��vQ�A��t�����Qm��+女z�ʱ�sM�t.첋_Ŕn����"�T� �@-��|�;����RD����jֿ�\�Q�{��-�{t�]��|9�[�9��l���AYC��-��,�S��K�l[BA+�e��*�pRٔ�tC���=�7�c���Ź�������dP���Hc]�˯��9ʎL�������Y|�*X���6��O�{\� CIM�,�8&�H�d�_/�����aL��,�=�� h�bw���H�N���4A���4�&$�Zq�v>��|�<�(mb=,��-�@���$�S���eı�n��=�S�'�� ���h�VE�dm<`��z#��]\�B˩g��Y�I��� Y�z6�D:L/��Ö�4>\ٗ� �-2���Gš�S�1�F/ԲTh8���l���T8��x
��~(�B\D~��hPa��|`�4�M�F����%�Z@�FF#�L�n������tV,��%�F2B��k�t����.F$.�+j�\Hʑq���c��ʌ�$��͝F��ÿS�, �$�@���������R�H�51!�tG�05W�	�^���Q9�A�/����,�)D#����4@�A`� ����U�r��z-�۵Nkh�t#	��2(����큌IZ�$���	�:�3(�@�m8v�ٮV��\_͇�N
���R����:Y͔�~���/��E��)Ǯ�0����K��q�2�S�P�������b�~��J�~�),:�����y�ۖ�x��M�:R-������ޓ)��Y�5�3P̿g��j<�z��a�o'�d���A/$Р����I�J9���p#0��#,�Qql�)f�>_�ܐ��q�����_�l��(#Y�*��I>#f�[gt�f�4T��pZ�`�ܴ��ti��XK�N�i�����Q�fw+7Fz����cZ4y!СwW2f[��EG��
�K6u|�م���c��L!$�v::�$o�Kiʁ�����ze%�p3C
sL蘽�a��"_�����e�#��<U���B(DQ�^5FnnlXd􆆃a@DX��i����0a+@��e��n#>��N�u����H*sGp�A��g�z��%
��rH�h�s�C��/��2, ��&[��1E(ߣ7h�/�D���}4�����/��鸂���?�[|
�*��OFeҧA�o�����H��͝	�pc�Ll�8�-(�<bi�W3#�"a��"a"�H��8ƽO��*j��v�r��!�b��T��)^:)���Ҁ�A��x��I�v�Sϗ��?��Q�Q~���َ�W�Y�$:B_7�X��
�VH�vl�&FO4��xG�j��P�Ĵ�ۯb��{��/
$�¼�4?�Zya���叼+.\��9��?T� y�4(�(9��q-��F2��,���ޢ��{�;-�V�,ZϮ,��v2��P7Z����D��0���~u�|�� $,:5�$p�m�'�"qj�&IS�� /�b臾�3e�����T��SΦBSjfv�"Ag+�N�d��@?Lۙf���[T�xV9��V�!F�s��q��9y�<�O�/�b�3Y^[ou7�1Τq�-`�U��q�=����r��$)�z�U�7Ƞޞف�Q���P.��&�]����t`� e�KVp� �͊8q.>�?d�ty��㋋�c̦��e���A���A���k���K�b��������>ܮg������z���~o��Fg����a3Q�漲�l���'=�'7Dh�7�L&���Ƒ�rƋ ��WO�5�(s��s����
��[=5��%�o���W]��ۑ��(�REE1U�-�K#@�L�k��h�X��fCK\���w���/����0�P����� ?Ü��\~?in%�& @�f?�$��%$ޥ��)
A�2��@��Zg�U�]��
��+�O��	�hI�x5��?���ZƄC�<�?�ܓw�̰�r��0E?�ւ�*
������^�edQ�K�.�d�Bn�#(���|q=������Q���M\�ƿ,�8h�'Ko`:Y.~/�S�< ����J���?vp����j��i�n� DhL=v��+��|,#��*/�Wf02	�;Z���_ ���F
1���n�g����4V�o���+�ԟDت_	
�G%,��8@P���i��ǆ#�L&�hv�z.�۞�`@WГ�E�$�	���G��[(��d�`oKF��&�\8�Ռ4�nc���3��B_i�%"��ʘ}p��/�vG�ٗ�P}��f\8�Q$g1��&#M?pv�yA�uq�]%����:Tַ,?J^vA�SM�3XP�3� �I-r puu�yb#��$gׇ��!�sg�w���"B�X��1�'���R�J/&(�w�G�1:\� $�2�T��G-��f]K���h�j�)���9�]MU~m�l�o�X���b+�v2������{��G��[�u��$tOwf��a���W1J �$f}�WGmX��B*X�/��p��W�Q}�m�1W��#�/����������I�!�:��]����It�?��Lgh`k�O���e����A B�f��*��M���k4�ĝ����1ߗ3A�{�c�Hb�_Ah�����d:H�� ���Ɨ�n;t�d��V6vP�8��ٟ(�d��坌4$��k1�/�����������bo�U�PcśdE3���8Y�ǆ![��5j�F�W���VӁ�&rנ�&1�[f���D�L��e~�]�t�����0��!E]�AÂ�JG4�-�.YApԺ�^�	H1�J�5��ۧ������J2�_��m�ƷMݚ$�Ȱн)�mǘ��g�7ŋ����a�i�!�}�zQ"!g�PcGt����
0�Ύ�^��4�4@��u+�I�^ƽ�?�A�+(��\jԁ���}0F@�
R"9�3R �Q�Ό��+�v&��hlw͙i-�RB���q�����B�z�3��'mH��n�6&=ڎ�l7):��6�ϿB�Aɍ��zV�ݨY�H͏���¡P�J 	y��9v���n�s*�s*����J-C�\"���cp3P;��+�A�4'�Mw��HjQά��v��*i��4H�:�(��a;s��iUZg�����W^��=}$
�1�ve�	8�戝 P��*�CF4O�	y���=�!W���m�a�I�i�U�R�[�,
�x;s�Nt�}S���)4,V�X4E�8 R�IS�z�!��%���8Jb�B�� ��+R���L�0�"��rr�5SO��Oa�m���Uϫ��И6k@};��D
���N�o�M�Wv
�"&Q8�Mɋ��YJ&X. {e�����U�~|�D�?@��`�/;Xd�[��#�Ō](���3�Q�p��n�}�^r����� P���u�ö�/���h]u�fd�M���e�N"
���+�UUy��c&_�4(H⩠��<�o&�B��1��A*
�z1�.4�A���,}ğAP(�ߝ��7�{�Q����:���=#�\�������|���P\q�Y�S��Z'ä�orW���S���/�F9�b<�5w�	��i�c�:~����4�/�E�� A�9R.�2���:8��XĊK�e��N�}�lo��H���r/���q��~{L
G���Xx��� ۗ@��<�/��
HXpt�������ntƨ�<�� �@�ڔ��M�#v�E�˗�q�� 3؁JXs�*���"&(�9��j�D�8���|���a��yj�Z�%��ǒ*�+Zjp?�{FP�<08,88��%��fMK䙞�+��,ǡ"K�,v��%O�4�%9R'���B��˸Q�lN���b�;����j�"U Ĭ.�F"����� ��@�g�X&D��͑�擾fm�0��\BQ7g��	c2cSJ?e� ��J���ܐ���6_!�L�(Ff��:�*��xb9��&n���W�2��K����F>��������CN���:�(
��R�P�%&���;M��w.5|pInNQ��
��:)QL��aA�9�vl�%C6hn�L��m�XT�n��X|^׎E�h����G�Ff,���Z+wj;���w���s�F_l�:2bƱ�;a�H��1�C+{�egG�|��1�����I���G1�we����oh��	^P@,y�3���a�RyH��8U]S��������H�X'�_JS�P�=���r��G��	י#tej���Ƕ���
MI�
�a �D��f�m1�$�:;�2鯸ӡ�8���>�5�y��`�Dh��ا�a�2�ap$B��B���;bR~@�c`[�M�Iܓ@���(��χ�b�pL�c��z;rJS�����#����:~rT�n����NC�`[��N<J73�u�5�r�B��-3�9\	��?��]����7�A�|��}��Hsg6�S���a@`UR˧��?�4L�lτԨù�m���WZ��X�;�;�-��W%k
���s�b�a�����4dXH�\/{a�?�Lꆉ6xw�Ċ�m&����V0h&��.��������$���G���lz�}W85�b[���+!0� cp$Q>���!h43;�F�~�|�fm�� �D�`D*;F�	��En v��������]���%��L���G;m�+���E0̯��yz^�������Ru`��%�Q�0d�5|&�U���[��qW���Z��������b�n����P����u{�F\��R �eP���L�%G3x����t�R4��iKH�H�MO ���[��> �?�1��I��7u���"�(�	��p�	SF&k�I3���:�<'ˑ���c����	BT�V͝ɏ���NQz4���\M��F6��+�:U�S��xBƌ�͙���8�	�?zλ4
ݬ�d[�r� �樿�>'�^�(8�ie�d�F���?�0���*�v�*��[86ddo�S�D��H��b�����sR����1B"ǘ�o���%8��ahʑ"�r��|�NLZIP�4���yj��5���13����f(��C�B*<���u���=�2/i��9�`x��t�v�2h�*��w��C�ͺ��y����_��-sy~10�Q%��V�&�j�oH�][�׈�����!b*1/��f���ċ�ئ%�&� �!._Gq=ԡCu�:{+��l��A�`Z��<zt����!>E1z��[�!�/�a�.	75�}�¡��Y�n���R	�'~4�|�)�#F�N(h&�ȅ�ar�NA�
��	� ��Ѧ�߽�0QBH,�m��5����B�E��O>P a��A��\�I���^=csw�ܟ~4l@3��'�x�p�Hܬ�&�����X�Em�kR�=�H�2|<Hx�m\�^hx�%]��d��������a\`t\����/!9n!w��_R:XS��wxL��\�N�/����/�B�	�artȤ����?�BL�m{w?�ʑdl�f�ё���ݠЪ�`���B��:.w�����
�"�:gQ���t�5M������Z%7���o�L���$�{�%4��M�	:��;f��v�	tٹm�	��z[cy
+��+�a��;�9z&�N�`�^<��RT7��|w�*;hF`��f�1|�TN��`��嚤&$Ed�{(tl����f�[���G_�<B��b��x���H�>�0�Q���Yg��!��X\�]n�s�/Oj��w�̳1*���ΰ{������[�}�*"3�^�3N� ������L"@A�L��E1Ł�dw[�'�~z�p�P=]�]��2Fg�F�Q��6g7�Y�N��/#�A*�MI-�2(~�M+攨��+�ceT8�ö�I������%��㇛����}xƲ6_}��(�����F��*V����ݑE.���W��<�-/> ���p�fP�[�O���ΰq7�� ��iwHR(ShbB8��I��py��R�_��I��aR̾D!;`�a�C�R���PK�|�\Ky��Αߜ����|,B��%
��G}��[N��S�@����vNe=|h���E�~b�ǃ*���`���S���|��@B���o���@=�}��5>�ZO�}��M�B�>��&jW��T߽�Ta���T�P�;u���u���q��f]�ۜ����B;��A���
(\*}6�����s�/��
�����UBG/c^˱���f;�^`?�S@J�ω������|&���4��BA���f,��c�"��Q����y�D�i�C%�������	��.������M���|�"J$)GSQ�Z�%���@e��]�L�vH��(��a,*G�����o��<�^U͝�jl��U̷��S"�������1��8M=�oԌT7*� .y���3S���f��Lk���]��R�������y�.��<]ͷ���(\wA�ˑ��������r�mB�3X�����Y|@��i(/t�Q�WI�g[M�b�	E	8��_�[��D�J����!FB�$2�r!��5܆���O�B躾�`���2�����)��	��~�X?ؐ�����3��	C�he6D����@ �ء�LǕ�T�
&̭���>�m4^��T6L�C=�`kݰW���c?�sC�p]I�����*x�����-7��g?s҉������	rs���Y�.?�AD�$3��*�(�cG����S����_ݻ��B�a&v�,9z�>���-�VAp~�d�����7�K+��j��nς�lm��H�ގ����ъ�,3�cR�T�|�����J��5Y	�ek���Ыe��W�f�㔽�P�\�ـ�vЭm�0\%���vLƴY�	�\,{f��Ei���BK��w־�l�K��`Pl�G�Ut��Z��K����?�e�V,><HW
`v,�4���!�G�3ۙXu�X,||�H����T�&�i���]�z��C˚)U�j�*ʍ���fBF�&���I�y"���N�]=�9p�Z|�d��j���UĖ�2�!��&�0�2��j��K����N9u�h� ���� nZ�rL$F��R2`5jn�?��!�����-�QY��"��C�����j�0���5��1��A��1F,p�4��Q���)�閟/�P|��	�V� �p�FJߺin�HK�w3~�S3 ��)A��G�d�����	~����򉫖����|�߄3Ja1��@�������g��B>J�ǅ�:Z>���܏�F���MGjɗ�����f�䯺^%y�a[��U��>�2�_�O\��Fh'(�A��k��+�1||��ƕ��\����o�{'&6�1A`��:Yr~8d&�~��*h�N#�\8�vD�Ε�޲W�֓AA�t��5��Y����4��͉��9�g��j�>���Y���� f��50�D��2�ط���8����N�Է��U02fI�������8�!���Um�R����Q�U��4�|hlp�JA�D�A�\%�-����A/gz��]G���� H)�^�rG�%�p�?��>��/K���_|�GOć������x��7L/���ea�$�윭f���~��i�pNn3b��Я22�D=+ō���+G�>\,���h�h"��s�u��_)��A����5��`;'�����/��P�H� 4p)��:Mԝ�Ʃ�|s�u�T���fS�00Q|����d���6���}�5��gW�T�&ۏ�S�AAB<�l�x#l����{M�Ԡ�I���
J\�Z#�&y`k�DfP��#��ص�;x ���6w;5P��qY���94����'���3Sx��{ϝ>	Y)D�>r
w���?�͌��m�~�Y��@X�s|�7�t�nF��߈�[o������F�0��J�n�IvZ�cC2K�P}�2�Z㱻����Vc�q���L�44Y�`�n���As"�@Ɯ^h<�f�?��-�?X�ʍJ��(�T �)%���"����IV̸�l[�؇����_eg�+���ݧF�[���&nA�����-�w�!/{�Qu��C���f#�d�Rok�10-�*���,Tv4�A�*r���1���W%z��	C��O�ثM/ʁI��T��y�$q���M(�j��Nm�3�NY�x���W0O�[�=(�����~�d���W�2�vߺ,�d ��9|X@�I
+�
�X=�;��(�)����w/��EAEV�4y���u$�6�q>�^��5 i�ِwal�PH
4xX�Pc6���!�z�B����;ŉ��_�1���v�b}�
Ж]��)�hD��_B��s����D����v�Gg�dT?p$�^é�B���n6���Z���逺��#��j;ܖ��=�S�'��_mZ��ζ�~�CF2�b���W @�da��{E��'i��Aa������|��X�����;k�'f���xd��j4�C:#kv`5�1�w®����$8A����'�y����YV/)����a�<nd��~�	������J�x����7k��c{��ktɚJ�o�w����rr�d9R�K�.�|!�:�S;(~;����&�sa���_�����m)i�@G�w������V����+���50!A��h�Y|DQ�HV�|X��%;	TяYn0�z���q� ��6�T�4���A�N_��b|d�(b��{q4����V�(�i�vƜ��,H;��+9d`�,�-�4h��� Qg����"�k�����S��*e	T�g�-h5@%C(<;���dK]0'�g�٬�1��-.�H�?��� A�G��r%�Q�n�>¥�@L���Y�H�V_dwg%672y��}�/��"b��o `5d����A�-���,u���Z�4@�k�F�����T�|�� D�q@����)d
+�B��@�"<��x��q��䉵�,��pD!��a��`��\��C[l1���A.1ݴ��8�$1����|)rY��f��g0��	�]�#K�&A����3���wpBa��K��N�q��y`�2m���
Xk��f���(6D	Ȃrå-T�#7��#�G$K��+�D�>	�4�vE�_M�������7�H�i
	1CR/eե���J��F�����$ލY�\�u8�l�<]��T�J�H�?��!�������6}�z��iV�U3�*|)��!Aږ�?z�w��5TouU�*9W%a �e�v��:n�q($����fZl_�j��"���m��v�ٹs��Ж�����zU�Q�j��)�ጾ4X���&0p�nE8Ą S0' -��o�����oz��kqd 1( �N���H��h]���4�ʈt�)��|�����-��,��Z��cBz����St��Ȁ!L�R&��/��NRs�z���G�b}�ԓ�Ө�B)��=(̈h�j��u�O�m������kH��$z�χ�:[@��U���}*�
h=�3$�>���>jt��/�Y���e�XUzY��1�;K_�E5Ґ���㸈��`I[sEL���MA����������
Eć�*��?nV_LID	&9�8M�Lk�4����d���i?\Bc�W)s�nZ}c��Q�<�{9(Q�;�R�@��}�u�
0ExH�����[��b���q��ʋ�1��1��%HZ����s��/�����d!�u��Zw���b8��O�Ҿ5:c����D-2�!��e����1.R��8Ҙ���F9PٞPT�D���K���.܂#�=w}D1��SO)�.��	"��㾗�h��J�Xҟ%���e��1��O�VrG$s�����/���I�D��ŉ���h��y.Q�}q��b@z
5
�sဃX�w��B50pu��� 9x�߱��i�<�Cq���ݲeVi��ߍ3�W�ya�#����@�"P����M��ū��$��w�
}�\�J-#�G-uއ�i�I'4���!�������H�a�Q�f��3��i�me� �Lh��(�74L �V��uE�*c�Mھ�������` O���#��i���:�Y�����X��>�)�����$�D61;tb� PI_yR��|��#����U!�%��.��Do��Y�
��1?qH*�4~����ɞ�S/�ӂ)dhs9$��ݲ��d4�Z޶34����&�,@������9r78��}1��3�-��@�z���|m��������r~�	�d�'�TD�_��wd%神�1�Fܱ�|��yH#V�-̞ 5����Ɲ��,���9����+/u���"ܱ�`�C	�����R��uW�[�ʿ�,�,�C�@���f�d��k5\p2���Y�HbFo�~s��.>��kث�ݶ�4�����"���Y��O)7&b!WS�|�8�T9���|�� �N(��I"?q����r���7��ku�o���M#�C
Gڻ}=XIb�Ԏ��RV�^�ljI�}���	h�x���G���Md��$N�h�
D�֫�N���F�4`�5���Q���t2�
�y�~5'�4E#,1�*!�U���V��3w��6QvPB-�1e��[��Pa4�p�M+�C_ʁ��B�.rMz��wg�A�&
�C�r�M�7F%PM����#y���#!��=�  ��l���oM�>���
N�eG_���+(�W�<l �WIA�e�G-��vS7�1�ۊ�%��k�s��VE*��H�H|�^:1(�`�]��S:AB�qtÌ����4�������JԎh�HJ�	��O��s/��$��L��|3ᾡm��!km8q7��%�)ڰ^t���-h�?.a Wͫ�Hs�C�X�t���N�KG���}G��Ɔ7�ٓ���PT"��&�ݶNX���l(�o���j�ն{a��g_��E��)��4�L�	���{�Z�Ƃ�F
R��K4��+�F?��e�$��(��D:��8e�u:JD�U���<ɭ�8Cw�x	g�0���_f�Y�Ñ��������q(��ů���;r�*# \h�&�ۆ*I2v��p��@dSa.�d3�N����}���"�O�U�x�L!춣3pܘ�K�����°������������e������b�&@F�w���j�����~�h��z˚I�^
�� �2%�'���h���?{��M����I(+��/�Y�� �bQ�Z���2&���?���0K}�/�Y��l��3��,m�U\���zue�v�.����m9}7pDJa�[:�'��G]��e�̸�z��>h��Ѻo�PA���	�b��+,�,��'>qu�+*ܵzS@�7;H�5���*M��e]�S��&W%���]r�8����ύvlǕ"fZ�T��RhЧw{���5���3�n�C:j����m�`ݶ��"�M���C���i��h�o,4y�ù�i�3�ˑG�K:c�H���X-'��Hԡ�=B�����8�:��66:�����	l�H��)������(�����z���uTk�Ѫ�+^փㄡ~��^��h��%���_mckj︒FZ��w��Īh�k��^_I�3�M|H���4=��D^�;��g�}k/��������j�&��$R�5�h�ń�^�w�7�q���y�?�d�Pr��܃,l�pJr��.����h�.��4�7wy�Lh>�,�#�
Pv�+X`�����m��]3o/9�� ��%Q��Gy8�h�|�G=*��*�U�O%q~��r,eE"�%��3Hg��UI�Li���Zϳ�0X/�v,@,�l��/'�C�����A�0
���W?��FGg
ʕ�T��#q`&m�$.tm��A��5b�a���6���|(A���
��N�:�'B��o��Z�澂ʂ��j��+�	0Ǩ���dA��N,�$��lju/�,�(�ܙ0�'9�YEa	���}�m�Zw�~��� t aB`�u���J�� �d�w�F�

:�w9�}AdH�İD+�P�|`&�,!\4=l�k�+�	����չDG�&|��|"6�t��u��ʳ;
 �S�`�.FE�[�^3�H����J/A�Hz��u��Vr9����c������h�\-��F�����q{�V����Rٌ_Cc�ß�$+[c�t�p�3"�e����C=M*rg�Qh���!M��O�G$�kx��qo)�S���q�!���B�02�]olȓf��IQ4}�9�t"���G���ξ
�1���]�����!V����{v����;�2�!#���S����"|�'��em界~������׉��Iàw[�|)im��A�K���_�wc�BGg��A��r�9)���/��$@����!r�Ev���ob�hb5�q��K�[&:Y�ݚdÿd;�'n���Ӏ�h�� �Y�:��7��ʋ	�o���+�h��h)�5n.m��U����S0L5۲�_tV�_���SY��,Xu����Ё

�(�h��ZH��>~X@fʏ}3M�|}ϳ}TA�S�e�K�	���~��n�M�2`ϙZc=��=����aQ�>�X��65F��}�W�_M����$?QWk���!It[�v9~������Q2�����adgi���"e�_��� �{">��4��d�P�[���=|<]P�ly��;z3����!��a�����E�o�$�kn�V���C]�qq, �G�<rz�g�L)�ˣ&�P��ܭu��6��|J��`�r)���1��۴0��lx�c|�C����c���ӡ*��<� \HhX�@�* ii��T�D����φ�Ӫ��PS�!b.T���a0Rb�~o�J��n�����c b��o�~�ͩ�k&T�(\<���tv�Ap�@T�$ǔ�(��Ai�	��4Fٝ���2
@��g���㒧�H����অ�_�#.s��ߢA�M&4�ݔ˴Q
�$�H����/ͥ�8H��V����sL;hEv��>m���|I>V�<����3�g1j��L��o��Y�{9���`V��-|%�jW��Q�6n(����3?+c��(Ɠ;��_�����'[+�#&N�v�B�_wܽ�щ����ݧoU�SahA�d���	���"V�
=�q�2�i�dIB�V�0��������_�4&�ĭ��%҃C+:���JБa./��� �����@����k�R)�+>C����$��[Ɍt���EN}`�ĵx�[�Y��p�4�q�a7����T,>.o��]�V��������G�03���9[���̈́�a�H�T���P\�>
�ѝ�f�M�'"����ҋ�B_Ïo�qз]����y��s�Ѳ�e��d%f�S�6���c�!H'�ɜI_n/-��=R�邞`A@��$T�r�Y~�H���(ҍq-]�_ ����D������`�+9(62Fqm�ňHiB�AD��o��r0��%��WnZt!8'w%pM���?�p͹~e������9CX�/�(���ad7����y-!6$�#����
XkQJ_M�d "lvyH�ɛ;x�M�i]�b~+�WB]������ز��!�;��E=,�0��F�@�IK�Ap���Ɲ\��`��G�
L��a��+|/�-�2a@f��p�����O@xZ�[(�F�N�G���f�����#C%�Cp!�{9�|W���7�
<d��z.�nf$�l�H������_�0R
3�ɀ#�	�X�Y�XM;�Sj�D���_��M��G���pLF�i:?|(�kѣ4�s�X:t�fL�j[M�H�� ����vL��!��O��ఫ&ܒD�Q�rE�"���"�	��jB����� ���i��9�����m�㭗���ڼ������%�1��,&|�w&;���*~4:4��m6�A��eKv�o��۷D{nGl���f+��
2�s|��^���Zn"�R��/�q�mY?�Z���	ͣ4Z�b�w�d���&�}��!�)���&��e؆DM��a��`�'��X�$i���U�7j�;�8��J���	N?*=�C���wz���é
��
=d��?l5���/Ӆ�kw�?p�9@��ށ��qRIq�i�<�Fp�l?f���ۧ^	�N���8�j��Ǒϗ�hn�Β@ӯs��)�,Ȳ��C}�%�wѰ�r�`�9��mq�m��*q�~2�U�B���p���5'��D\8�[�Ja�#x���m�́YN~�%8��x�A��D4���e���|�i<q;' ���F|�֤�&��w�e�&���!!tƣ�9�/�B�L��5_\}Z�1�l�������T��P��Lq��8G���.�;&␳Ȗ^+���1s�������6�仡����*�ڳ%9�ʹܨ�);�����<�kn��L@�/��<sN�V)|	Z?D��{�
�ؚ��1�E%���£d���}� $@�[>��0�@�������CƇ��uB�h.Э�z]?y0��v��1_LYE�_�ƄJ<�"Ew��r�~u/���'Ff2�("D�=l�w�d=;�4����g AhQ�?��|��V�H������)�&�_$���$��p�CK���֐u�?��7�R�r�8q��l.Ñ�z��;��,f&R
�O�@gB�&�����&nC1&N�'Yd>q`�:�&���ln��S��.�����U+�@�6�>�\X�V ?�o�\f�
���R\��&���n>�m�_|��SQ2:/[���"++�����w�tٖ;BXݽ�x4?��۱�z��+��,8a�[��i�1c~�*e�
���h�2�v4�c�.�5G[�q??aЯMk��4|Y�����k[�/>��tmg�b�\��uݪ�(�����0*�������B�Ǭ�GCщ�o
Fn�^,��5��b	Yr�W��
�@R-��1�� ��G��"���a�����m�Z��Ieb>t���2P\�\��Ng%�0�G�x�F���k*��|�=��/�b_�@��Z�67��k�[�}�����@�Фb���=�b���@�F&�[:����Ղ�.7�����~��}�e�+j���DߌП�!��_m�6�f ´�E�b���E����)I����+�=��:O�B�����d.�F���Ӷ����P��$0��m6��Q��1�
�Ԩ:y�u�El�C�|���7��Z�1��}4Da�(L��ih����/�F��!S�]���G9/�A�C����e�F(,���F}�#b�?�(�����x��8�cqg�D�	��XuK��nV2�k)}�-��C��Y3q\}�LR��Z���J���A�@����rC����t��d�	���)��t�����������Rۓ��)}�����eb��o���0�yy�]4��еM0��&�y9N5�ߦ0���J�1�=��^.�z���0�^ۖ]K�v]i�j���3ZC_������x+'u�i��0�L5/���!�3��.?��H���W	di���̜��D1R���r�H1����	�h��m&�RZ�|-����D�?�⡭���A���ċq��5��1ߡ���da��@b4�sh&
Δ^�#k|��'���O�c&�zRk��/���q��{��ǲ����}���2�c��G���7�r���!vNv�o��=��7FLl��[?�iVw��_���i��a���D�Pʧ�|�L�p��["�F���{��v.5,�[�fEU��Ft�Fz��D
�\5����}�o`!�H�x����e�N��fn15fCB�i���%TZ�b��2i܉�D:�s]���3-
spF��7H�w�)��hd5��70E�1��ŗ�k�i؂�QFnE-ehH1(#]0	},�"]�A�yz��yb�VE�L=.cEV@sk�'���ūi�k��F9/�f(La#���e���CB�����
�ٶ�(��Lm��8�Y������|[�������Xv��2߹D=|/&{噰�+�%6��6s�|��z87����D;	�=���8Q�t��,\q��Q��!&�͟�	�0׻���*8��[[F�B ���~	Q 03r��bˆ����w�PxK�w=,	��#��9�]���1�i|��ZA��wM��Ȓ,�i}������g�6e�QܾB�I ���~X�o3˽qlۖ|�d�_0�d��6l�Nh��	M�aA'�;�|�Ӆ��	V���Q~Wa���+8R{�7n�`ϘB6m��/��.,H���d������|�E�se�'�H��}�r���+��Cm2	8%!*V�g��gQ��y/9�A�+6���;�B��b�Ds���M>4���q ��w���cѽ�ѡ���R�Uㄟ��4kԕŘ<s]��E�Ɓ���ײ*=1�;N�nύ�wF��*��;�F�vqi��&���˽��[������Ļe�?_�f���aA��]�fj�_�5>^���6N���*q�����sx.H�����z�_�.Th"��~���O�jm`�sC��U����)[�N��Y,�9�~ٮ ��)���K.�	'�(�*�g��$r���ɓ�Ƃ��[��'�e;ٛ;�I��:,=�^�>>_��Pg�|���@��@@�eE�Q9��ż}�ja}�Y~���aS�+	��ֲ�W�PL���l�5&̕�f0�̸�m�~_rJ%�J"(Τke������I^���j�@F����ć�����M���	[���+)BL.�W�;�ȃ%�Qw��7Q�+č�>�
��7�� ß���X\���4dj��;<kD3�D��6<�IVx-�_"N�rg�5C��Ւ���<������!�����b�O�r~_��S�.��AF�Ce�v��\�r��?pJv�:8�����}�N���*��o��A���������a�NE��\-i��@�X=�A��q�s�E�K4
���Ow5O��"m��A�VXT!�џ�R+a"�[<�����ė�g���FZl!^�����D
�i��p��B�!�m�b:/,=χ(}��n��y�ݺ�a�n��X��xQ���[��i���%^��`�XC��#n~�UpM!�i/��DJ�k���7)�#%٤Ðzn�`�f������| �nrE3,(�[t��!$�=�	�1���h��z��-��b�p�Y���|�cl��!m�/_�TIn�n���Hv�ץ�S��Q&Xb���MyR����#m���)XC�!6��>��J~��
0;���¢${�p��ni�O�,�����V<����<O/f�2�`�Sd)������p��y"ӯ'D�H���h"�/�[VA��4Ycf ^�ɐ��`y�O�{�Ď(�AT�(���/����"���82�ӉN�#����%��mE��'Ec�$I@wN��r�}l�<���D	\��z��V�| ��d�@�2���X�s�Z��Ӯm��1��O���wq���]�R�����Rb�Y�@��0�Ev�!��U5 " he����6?_m <���C% �ߪ�C���H��'Ɛʧzh��c)�c�i<�y��O�Z�9s;��!����F<`�-����!8��z
\V|�>����~{$��"�"{�~�۲�����c	O������><�\U����IN(�W^L��d�r�.�a��m>کe�&E��n>2��*�H�f��*��w5��Y��� �O\j� O���>&/h\#x&�$�#�z*OJ�t����]���\���za�
��e���(V�M9����tm�|���Ehtb��4Ȅ%�Ȱ��c橴�d�֕NTeo|Y
��~4q�zi�􋛸q(^	���D9A��ݔ�Λ�7h��4�A�/i�{rs��	���%���]��N�[��oE.5LgG�0+�$��/�z�џ�#9#��ٶ�G� �^<m��1.���WB1|ŶZ5�����Y�r�?�s�#jL�n���ؕ��Sַb�r�,_���.#C�b-�A��9
����@AS��"�C���wm��&����n��Z��9���Ң�S�87�����KF�&6[A-��?S�f�<M�]Au�z�h�-�L8�<�z<%j �������{%���f�M9!�;g<`��m)�Exx!9H�k��F$f�o�[��^�F����1��F�&�eO��\��=�χ��߷O�*�콨&:!j˻'�_��	�'�1��L�&��ֻ*����X�Og��
�T�t��	���G>	�h�Ϲ�����S�W6���d��L�/�-��-��<�k���V<ĠD�r��>_Cr�Ru��"��~2������ǠB@G�m�[������ye`��R�@��	B�m���ۺ�2	p9�7"�����ɘ7����KG�}.̸�
��^2�U�X&��q�vN|�Y�i&�e33�v�	
@A!�g�8�G���y���ǎzo-��W��,��ўi��Ci�ϔ��~
3��T���������h�)	%i��N��8�c�9�?�D�*[�����)�so�K���� Ҡ��J�";�y���{���	�ژN\�α�Y�]j���g�Jlm���pU�<'ˏ���e�~L$���?S�GBT4�
���TIWځnB��Oา��%��§.}Ӷr��Q���y3=7����	mQ�[�e��㏱����:�b-�s�=��D(t�Ai�t�[H��Du�4Q��n�#=��䆚��}�J��)�f|��H�*���#`�6��r��'W�O<��$"e���-Zv�!;6s�]銛�G�ţ�7
%���g-�ab/����Ӊ��#&n��_h��I��w�@���)�|?�1�ѷ"��x&(��
�y#��B9h��c+Mrx?62(\AP#I75��vIQ5wE�|*������l��s<Xe��K�W*m"�H*��/��S[x���e��	�]F�7M)ʸ�nbm�_ᴝ�4.Js��f�u����|�*��@�@h�v��a�{�VL�5#�CGN����_푤#/�D���Бy|H�ȁY]�M�,��o�Q��eM#��g�!����Rρ�!���8�d��(���E�����N:l��!�B�
�7"�ՠ��[�7n�l�qX�NP@K�1<!�f;��9dm|���05"���)��/�R
�F�_�DS��*��#4LI ��h��Y��ƂJ�ߠBG����f����o])}�		�C��$%�����z2�o_ݶ�˒����q�0�,F�B�EGVx5��ql��J�����3���i�.�0A��!2Y����?ʌc��>_9%0L%�2��#c��!A�/��cKv�8�$i�{"ќCq����^3�y;����A���]t����/�*�H	���e��Z�b��}eAB���i�� 7L��-Ӯ�!�E7|B��U	��D�
r'�1�)�M42�2O���D�۱�2�@&:����ﻡ{���ov^D���h����#��7h�JF�g�s2�I��]��Z4�����Jt�;�=g9��E:R�'~�@GK���>j�ho-��D��kJp���q�WA��S�9���J��hc[�!n7�k|@�	q���pB4�U��q\�%�V��A�6q�*��k���A��zH�K�P�<cwcs<�L������qV�&=Gr��[�����¹�sL;[��|+��V��O9�]ڽ+;G:ə�|�D�y@C���۴�܉'�"�	�<��w=���S>'��˨�H��/A���3�����wW��U`�����������m�A1���X"Ը��1�g�U�D-nZ?��<w+�~G�ܖ��ϗ��|�ec�$����f�;).l�v%��
�&��|���g��A�X%x�V�g��D�@T/��Hm���`Ѡg˯�YE�d�	��������Z2+��6�*5�cմ��;r�G�3W�ROr��`��@.�I���
N\w��=L��PzW����C+�dxΝ��_������;�Z{jH�5hQQd(���<g�����|�G_,�d�s��,s�6~
����&H�ȿ����	����h��.JW/��X�:� a❑�/ٮ

+��ws�X��c��QP,	�Y�@N�����Zsm2�-��؊���,7�ܹ�����V��a:��'��\|�ϏQ��Q�;�"F���1q�g��Xٲ�M�	.;D
7zF�x#�<���Z����>���L��"�;�f��)���?=]N;鳰D���c���C����a����止����TU������O_�(�G�Ak@��L�?�4���*k���{^�٩س���%%$ʍ���o�������m(4�s�>R��v�mXM����7h�Bcw{�pBB���𠓤x�xr�4]����^��q
��X��rTj��5w��`.r�N�姿�~���;�Q�%_iڹ�lӮ!3L�����&��
4�3��Fv��U��h�[2��َ܋|#=��c�A���I2w,#%����x-�%���{kK������~)0y�6�+��H�"�
6k��˱����5�~0��Zv7)PX��\��)=f�����N�x{�����ȧBV&�� �ie�宨�PQ�Nt��e-���`�@��[���k��.Xq�roP?�BAέB5���Xpë�2��*$D���6^V󽇡�|w�pLd6�)�U��.x�.����1[��児��&)ٌd��|�;�D~O���/�K�=�힖�c��Ph�A�?wA)ai�
!�Q���Z�v"�ǜ��߂S$���i=낱���4g��ml���V�w���+1���Bͯ���¥�r�2��߂Tמ�ߊ��]�����C�!���S!J$kFSe��r�Q�=<:9I�۔ki�d�ԻO�AC��iχ����[f����JZsaM͔�scEQo �Wإ
W�AWs�w���G����ݤ�y)jV�.n��S��	����y�_�'��I�����m&>o�ⱏ�u/������1wp>�8�
E�h�R0Ec�,C�ſ�Ǧ|rۉ.m�-�⑌ɷ��%���mD�}�^��J������"ѹX\F�^�x'�7>+C�"�l��3t��I{�&�7F���=i�bT�,���1��z�^	q��A:)hsV��)�{बc�Ã-��=�C���{n+���7���ރ��O�av����Ħo�q�Z{�9hȾ��.)I[. ����BNAn��[e�%m�@�>	��r���$�S~������x^�M�h��h&n��V���A]����.+��"��U�| �����Ad$��MBR>w�%17�S4�F�&9����o�D/�߸+9��E|�,*�����-�s���8����3Eso|�ː��ٯ�L>��&WHi��[��qi�=�h�>�$q�)PQӭ�1m �45T��c��H��z2i�����<>C1��/�W�

�s)��O�eN��R��;��HY���O�D$�4��]��d���b�E�^^����
�wn�8�t��h9�Y����d|�\�N:9H����HJ k��IQ�'E�Q�}�鎜'1��W��*�b���k0� $�	Q>�evg��A�7��Y�m�FFXf:�pHJmʺ�𓏴q��
}��@�B����A�>:>�wm��E�E�4�ͻL��r��{(C�c`gJS�G�<3����w�X�QR駿�VQ]�<߉�F8׻�%�,)s#��3����W!�~�7�e�՚�;v�I��#sq/��c\H��!�ŵ�~�0���!�+ur�c/F��5�|+��Q��K��۹����TZ?1����vv����%Gu��=.џ�@ix$SPo��]�Wԑr��-�y`x���I�p�ę��ਆ`�y`߈}���_
	
�m{Xo���ҫtfm¿�'���w�Jko��λ�N]��ؤ.VH��G5�t{�7��;'�o���I+��`p;��6j�?����x�����_�G�{�ǻ�)��8��=��i��WJ�  ��a� �_ ��� ����ҩPƼG֢�6�:�f7�B��@���<�_$�|G#6��MNw�yJ:������g�TF�MYߝuj��^	������#������R��+��!�Zm�A�U�i��[��vݳ2��aJ.B�O0[�N�pe�H�A>���g2`�Ƈ��AW�jd}��y�,�9��"�x�� {̆�o�̔���lm'|?{3�M1� ��q���\:XA�x�m���|;�c�*wK��	�!{:u�������Q�l�j6͸� ��t
��?�.�-�wk7_�Kh��硵|偤̤�����xH�j��*%��1�u���1�� !g����J�+4O����ܥ�j�����K�+/-�XW:i���!�5�3=����NI�`Y_���{�W�i��#j���B����_GhK����W���ص��c��}���&�9�޼���z���bv���$6�`���TP������E�;�������۠���P�=�~j�-�z?	c�/�ݏ��n�}�y�%ڵxc¤��i����A�	�K�3��n�|>V�-��W}��hg��o����-8��a�Tt^��RX�[����q������`�Z�Z��Γ
(ٹm�]����W���r�e	T�?4_m�B�H�G�D�X$GP��&�.��2e]/��t�B���}�1�d�z�wk���a��-i.t���Ѱ��n�