E�j�9�,���U5ִ��d�g��Oe���L24�-��*]�&_�0�H⻰�g�%�D�y|����l��H]	hwBY5��>�n)B��^�V|�B
�EaR쒾L��5�I�aZh�v͡7'�#���Y}P���`G|�4,j$�UX�_%�`���V$D�/�m����������\xMOVH5J�(3�5��j�x_$�P`R�C.w�F��� R�mA�Oe�Q"L�:9|Jq6�����L-6��J���lH�J��8�:�1dm��eAA��I����_!˄�����T�|M��y�@]�"��Zz�%�S<�^�`�Fׁ��A] ����l>�2K�I����*�H*�D�͠n]{L��3
�y�qs���kw1�v �h,�r㿉~[Hp`
�w ��7����4�[�����$ˎs���%�W���PN��������
I�I��
���/��X"$XL�8ޗf�"��Y"�� ���+���)�CSQY��;���Bm#�Ơ	�_��ubJkH�X��S9�TR DӁ�i��ŗ��(`'P�G�:�a�_?݈����Րo��_Q'�'�>+�ة�ǌ�,�W�"VM;�A
]�Ju�J$���"��� T�t҉�tGc�r�0IB��h�̾!�#�G�$P�+�K���\VD.�_A624HxY��%��
E<�NiE�lC�E�L�u5�x��������s�gÊ4��>l�q���\f��P@@	aB8�B�I��T�EŶ� ����_� *1(&F����6��K��<q�+B������	P��(�{���R�[�}bĔ#04.`�P�-�#� ��ϫY��|ղD�K��w+orSd��d�J���dGlHD � �A����bD�%�ߗƍ	!d��%�iR0@`�4�V��#���P��ԆJ�-���\�gS3�р���
��y�u0w*k�$֡5��6Qw��D�2�֩��� �61zJӇ�������P"@�H�GQ�6�jfW��"$k!�Wq�J��v�6"�lYVx�lj_$, �.��V	�ë��-2R%� ��w{
 Q1���*+~�4�R(�v�	"$���n�_�+��a�K����Y���u͖�%1�V�Ĺ���zͦ9L�+9��%a��3��"H>�B��N�qCV�vRl�r�H"-�5�������Ti39�ń�j�z��@ȰE�K94�;�		A�J!;G�D�ܸ<'"D�|t@���5�p��DQc��/�AX�FY���0L�8I�3�z���Dq�P�%����<J��"<��3�/#��y���K^,�<DbĸH��e[f��7U6�TT��8Ҝ�g�j�1�7e�%FP����������CY�}U#U#�~�I��t�����Ae�t;��.a��&�a����`}�~k�$����<�yF�F��Ad�o�j�9�3 �]��5�xdV���/��,$(>��\>I*�f�L���(���Z������)x�������~B�<++e�Z����x��
 @+Gzj̿�_-��%�
Q"�7�x�zNC�a{��m� � ��/��Kȑ���U��k4��W�3��w�G�cJ|-�X�ylr�lQ��9����p�H��(�a�������5E�n��4��d��,��_AC�H:"�(��G��*J
��G2l��4�4Vm��ܾ�*:F������_apf�(-����
�,4��ZR�ЭJ����,m�4�i�	��3��Xȸ��kҺr��	��$� �,>�q��"���<>�wkVx��`��?/� FAL@l�B.Xّf!ΥƸ�UPm���� `��+�lqB⿪�P�d,�(X��5��С���K�g�uj�@|��	����.W�һr�cA�\M�e��[�PZ(�w�K�8D���Q>��ͧB_
�
BL$ Q�l��_����q�#�w�((���������պ�/�8D�l٘��2��HT+S�sݵ��q�tC�kwv�4K�-�ޯ�2�U}fS����Q�1����}��^/P�����dY���W��3��"��V��Vuf��3'hG[N�^�0��jK�4-��E�^!�Vg��	PV
M:���q_$��Q@"�@�m�U��XQZp����n���Y;J`�k8H��eNX=2��|(�ja}�;q���$����k�ŕ�TWOq��Y�d��L��K��R!6B��B���>~�J�/��\,Q ��nIe���Oq�$<�.9�[�Ge�����-�k�!ؐ]>���+�/�HQ�$N_�CF3G*��C����V��(�LRb���|�1��(,- PT����q+��Ņ4~Fnf��3(�s!g��$����аSx{8�)���>"j�esj�;\���$+#��(�g�twx蔠��ǖ��w����\����{�Ȩ�J�K���Y��C~<0�oU���Zʼ|g�UZp����w�t��{�"T;�ډK���N�%�/�[#O�YiF5Trm�!��bxf�OΏ�E͈��@e��M��w�R*�$j�~�0�=�t�:nP� i��b'Sh;��
��'gm�#�T���Y_��& ���rܽ�R�)�;�����-8��+�B8�����J�n|�|s��ZX�H�"B&�T��s�e��$@�o.)7j��;�`%��Ј�i�5J|��,AE�z��&�w�E�S�/�)	����mGt!���z_� L�YCEܓ_��đݒ	Ie��
PPX=�j�m<e�����6sP�G�fW�:O���9|ѡ���Ta~� ��ř��9C����1���N�D}:^�`P�g�\�|H��H\bZO�[���wF+�v��
!#����V�MF[�x*�1L��7�w��䰪�s��d8/���Q�[f勶4��cAIJ?��Xl*,�	
	-���B�Ҫ�m�?�����6%���p�ݶ��f�X\�����*�����z�����/��XXPD��ͦB�:.L��CL���me�i��ҩ�L ��M��qޙ-`w���fDL��Ͳ��!0�G/��Q;niQ
��$\�?J_$H�B��T�O_	��*�n$O��r���\���
ŗ�
8lH!n]#�;cr+���>�F9ѽp�Wf�2��|�k��RS���LfM]����BF�5��s��l� ���^�3Q`Dr!b`��(�iQ��t�
\����NND)̃����ω�.T]�T�@^,C�]��v!8�x�m5/���&
�D����~s��S��x��.���p*�j!��]F��H_`*8LaB^��!Ø;خ��L�F�ϚE�����[��r_#X�!���H��$�9Ha��$�0y�-��,�	a� �[�����銾	Jl�6����Jt��ғ��v?"���	]ޜ(�^Q�\*7��Ĭ���0�P~��"�c��}v(I�Ʃ$�Ё�ha���¡1+��4X"���p(V����܋탁��A!��Ja�'l]r(᱆4��i�&��n�w��F=����K.�1ߤ/���)��dl�w��(��@G�kv�3�ܒ�7�@ڟREc�k[-�n�dKn�Hr��F?�4L8?�@��Hȥ@2J�8v��D��ި�gnW�����-�Z�6��u^iD�L��gt�.�ˍ5N�pĵ��������/j�
�Y����"���Ț����
]��;e������:I6[~,�^3M#V�1)�i��,�_�$�f[V�ũ�x��,<e��ǋh���3x��Q{��?e7?~v�rO�#Iw�&�*�T�AI6���I'ˍ>�?�����,�(�Da=ˉ3�َ��j>%�*f, ��)����g<d�e��D�)G
����4P�&M����1��+������[��6��;���Λ��ZN���e\WbC�B�t��Oȋ��ą�A#����e�����iB$⹡�1����vM���O��r���Y�b:������� ���V,<B*��Y��ĜVT��� �V�	�Vn~�w:�T�)�i� �	�o�8�zy�/>f�|;!�8��Y_��;��4�l�W���C��<�g��.�^we���n�� 8�/)`��حo��������dKX��С��HPL�@��4ԻD��AbW50�W�Q托�]2��Y�J_(|xLH�0b?��7�'Ƀ�]�Z0t
@�aB�;Gp���8Gc������'��d�����yΏX%��|$-�(F
>$�!����7k�|ef)^�f�fl�udO&r/�'i?��H8<(�|�f�yX�]UJ��tQ[f�[vUq[L��e��	�0�����\�Vw(*�H#��Z���Jcr�t���[ݍz��W�S�8��D~_�^�SP;�NW�i�~Ŕ$4@�RA��M��l�8��a��}����g�o|�6�db
�yJ�1e��Ƀ����A%wj�j0�(�V�'����*���U��1^�K��x��j�4*����z����-�^!��ۦ�2�����͍�� �Q{(Y�!{r�X�S� 'K��Yg��$" x@ R	�;b���cE��4��Vڿ��%�'��X��+���b��)/��_��7���d��D_/��$!B�
\CG�\?�&�����h>t'ZE�>��!ANkܾ,����lݼ�7�wc���Q�h��\p��$�pʤ�ř�L8��u�鈉ݐ�\��E�)a��%L�U�{�''	e��pr��j�k��6c�f�lV��FߗT� �����ca���b�h�E:����ٌ�K����a.9�h����ɿ�k��DG4��/Іb��u����]�;�B�N3��V|<�����;6�m�i���1�I.s��R";`�Hf�Uc�.'��~=���&�٢0e�2i��z&��eu���K��0���	�%�(L�b6�)2ٞ0͝T�c_niJ�ŗ����G3S�O�b3R�y���,�J��Ih���JC���֬������9���F�fl�&K$`�{�j��N��j<X���+2M���=��Ǯ�4`dP��d��7�'��	�,mKY>�֚���B�	9h�s�r�Wtc*��o�Ln_G��_m�0���*�.��x�J�@��aA�1��;���'���n�*�v�͙��!ʼ�+ж
��Fv�&\?S|�	lӃo�sz���?˴��(P�I�Ĺ>E��|���O �
K먷KhV-&�P�{e��,HKM�V���)u�.�pF Q��a�8�>� �A�~�3��e� l	!�I��ze��LG��R�*A�Ͱ���O��5���`ɠ��b t�u���а=�"`�F;ìؔMr�����iA�z��{Ж��\��0tv�Ժh~Y?���/�(��H( 8�,c�.w��%�cl�9Ó{j*�U_2Ԫ]a�B
�����h۠'3�C����
���
	�����K67+~M6�������hXH&9p���sw�0�����7�9��t�ʥ ���nͷ�[31Y�O��G�e�T�fm:�'���l�"��pJ��0��4�B��ʗ����I�����V�.sxj�l���v�</V���yx���S��|��
*�~s+?���^_/�0B���9�Z��v�_�8������e�H A��YT(�U+\cC�Ɯ:����3w���s�(���^/��," @�L-=���iv�لc���p-r�.9�t8��ݹsp�*���p���"�������H(���pV�^�u�1�Kwf�����
��V��� ������Ae
8��:����e3����.>���F_^؈��L( xzX8VݠH0h`S�P�R������O0VJ�vY��0v���N���� (Ml�kb����w�TNM�L�
@���»\L�����q
eKLrf�P�n�6U��w�B_�o�����6\4��k,<L6�4r�j�M/������^���I�-�(�����!D���F�y]�#J�.�цVu�{�Z+Q�R�r�#��M��~T�n>�R�e��!��i��FӒ� �5��h�q�l������!͐����r\/	��&^̷�,]�/�b��$�[��Z2F�Z ����ޘk�Ż���7�7�.B�V�7i6c>F(`�Qq~�J¡@��>�a�q<�c/�}��0!}���NбG��M��X���,��]��_D	���5.���,X$y�@XA>��1����2�1fؤp��� z�s�`�I^��_��F#\�>E���65��|L (��F	X�,�	��
�JMȰ�a��w&t{��!Un�V}��FƤ�/e�� ��('9��닖��1���F:	З�.�L:e��
�@��a�1���?*��P�|6����Q��&$�L(O��G7 3��ٍLF�ձ��mϞ�V��x�+�|	� Q�\�Z�갌�[l�B��S�(�yy�x��
�D0����t,�{��<�b�[��8(#(�I �*�,b	@,�<��
�F<�e9����w���r�q��u��狀����ロ/?oT�4��U�qF��mI|0T@�vG��@5���G��aUQ֑*�����.�9I���#��#ܽ���;�n�)fh�x���D������� �\�O��e�D<�� ���(ΰ��CG�`�U���(*
���`�Þ��|I�"$}�<�\L��S��*wj�,.V���w<�,�P�<�¤���ﭞ䫗� �8��'i\��~��2����Htqx�r$l��]��O�	��T&����mt�8����0��$b�uI�N䢺 T=����,s��a�`{ܷ˄�CI������LX�4�]"�����2MQw��ޯ�{(���B*A�ipX��3��J����r�\Q��'�ЁB��,8�_&)���/��	PA\�|�ѻ�4���"�2G��cO�_� �Ә$$c>���o�3��2�W�F�UMj�H.�'^�b`_�l�R�  Á���B��a1�Ш<��8��-.��XD"V{R�0ú�' � ����b��?�����.����O3�w/:l8�2�K��<�X�����������1���iP�L�#<��(b���C�M���q�z�M������S�G��ە��G�$�H�~�xƯ���G3S�j���Nx<X֚�aӎ��^[ځ:#�W9qM���j��ȋ_�- ��N���3��ˤ�Y�j>���$Zi��FD���~��0;I�3�����>�6��A?����4�?��	5_v��eTN�Z��)����'g4ۢ�:��HE���r�1"���
G|9����c� vA���b��E���3q[���"-B�9ԕm+����"��� A@CRU�{��(�f-�/h*4*� �ٱ]qj2�˗9�#���S�q�h̑Ǜ���"���p�6 v0	cN�˂��'�y]��=�ɀ����4ߗa\+ɥ�v{2X��s� �ÈC���Tx�k/�	����0Q�9n�<�� �!y�F#��;�f@~J�|�c�8���_�䙙�t��ȫh����� !KrcŞ'B�a/!�3�lVj؊��̾�A�����0�9���g~���ǲ�c�z�}'��[M8�v��|5���q�"$yM���K���p�Y�!�1e����p��c��L�R�M`���=�ɹv6s/��ㅂ�j2�b1��6�@��Kc�w���G��";�Ƅ>�\q]�p�D��I�b�]e�T��0���,gp�t@B f0����B���
�|,r�\82�ᣒw%�k���l�?��
	'���$�,`D�I��'��yc����JU�>�[���B	�?��`@:<i�'�/'�D�A�QO��>|1.2H�hp���&���.��{���$� r<{3B<�c/�� � @�+!�Tܷz�fS��`��`Q���ݦW�}�� {���$C�8��|��"+�@ܐ ��s��˲��E�0$0b��,K�4��������)���^j����EE.��L�oS1=��	�RU�8�6JW�e5�u�ɽ.�{��v()Ӓ�<�j^�G�_a"aB�Y��}���iH9$�;V�����UD�]�$4@G*D룟F��.������B�ԔR����a&!�l����q��tQy`S��^�#5̓&e��Nh0t�"�vL��2B� �E�f�BX��]ӵ0�dcR�`��Ko�6~{1�(I��	V�>P�s���@{��I0��|^ݷ.&iF��!�\8�VQ_4�nN�|�W�l���]~&������G�jҩ#r��>�C%|nu�v֏��e��1���l�;N7�|~C*�7��xH�\|�u>����d̴K��ŐDt�h���=5v�yB'���J�-�r�����6��մ����H˦����t���.i��ѓ�%qU/��6���c�sr[1�1�ě���^/�l��"g�>��;��2(�������!Z�>�!�*�}D��	I^ܻ��`z�L1�'��9�(�[�/�$�(%�dl�{��e�A�ѡA"Q�67�� �
�lPO���_ ��,Q:�/�d��6`�d5�K7U��}>�H� z�V��L� �;u������� �ʪ9�$�pj
u����\b��P�e��IJ@ �R�%�M�o�_���]VY��E��;�Ѡ�0�d�v�l��1���XdN���ĂL"@�Ta����q�K��Q����XdH-�r5
�"�FV!eŬ�82C��#YsVf�b蛜o7�f���s